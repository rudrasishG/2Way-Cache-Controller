* NGSPICE file created from cache_controller.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

.subckt cache_controller VGND VPWR clk cpu_addr[0] cpu_addr[10] cpu_addr[11] cpu_addr[12]
+ cpu_addr[13] cpu_addr[14] cpu_addr[15] cpu_addr[16] cpu_addr[17] cpu_addr[18] cpu_addr[19]
+ cpu_addr[1] cpu_addr[20] cpu_addr[21] cpu_addr[22] cpu_addr[23] cpu_addr[24] cpu_addr[25]
+ cpu_addr[26] cpu_addr[27] cpu_addr[28] cpu_addr[29] cpu_addr[2] cpu_addr[30] cpu_addr[31]
+ cpu_addr[3] cpu_addr[4] cpu_addr[5] cpu_addr[6] cpu_addr[7] cpu_addr[8] cpu_addr[9]
+ cpu_rdata[0] cpu_rdata[10] cpu_rdata[11] cpu_rdata[12] cpu_rdata[13] cpu_rdata[14]
+ cpu_rdata[15] cpu_rdata[16] cpu_rdata[17] cpu_rdata[18] cpu_rdata[19] cpu_rdata[1]
+ cpu_rdata[20] cpu_rdata[21] cpu_rdata[22] cpu_rdata[23] cpu_rdata[24] cpu_rdata[25]
+ cpu_rdata[26] cpu_rdata[27] cpu_rdata[28] cpu_rdata[29] cpu_rdata[2] cpu_rdata[30]
+ cpu_rdata[31] cpu_rdata[32] cpu_rdata[33] cpu_rdata[34] cpu_rdata[35] cpu_rdata[36]
+ cpu_rdata[37] cpu_rdata[38] cpu_rdata[39] cpu_rdata[3] cpu_rdata[40] cpu_rdata[41]
+ cpu_rdata[42] cpu_rdata[43] cpu_rdata[44] cpu_rdata[45] cpu_rdata[46] cpu_rdata[47]
+ cpu_rdata[48] cpu_rdata[49] cpu_rdata[4] cpu_rdata[50] cpu_rdata[51] cpu_rdata[52]
+ cpu_rdata[53] cpu_rdata[54] cpu_rdata[55] cpu_rdata[56] cpu_rdata[57] cpu_rdata[58]
+ cpu_rdata[59] cpu_rdata[5] cpu_rdata[60] cpu_rdata[61] cpu_rdata[62] cpu_rdata[63]
+ cpu_rdata[6] cpu_rdata[7] cpu_rdata[8] cpu_rdata[9] cpu_read cpu_ready cpu_wdata[0]
+ cpu_wdata[10] cpu_wdata[11] cpu_wdata[12] cpu_wdata[13] cpu_wdata[14] cpu_wdata[15]
+ cpu_wdata[16] cpu_wdata[17] cpu_wdata[18] cpu_wdata[19] cpu_wdata[1] cpu_wdata[20]
+ cpu_wdata[21] cpu_wdata[22] cpu_wdata[23] cpu_wdata[24] cpu_wdata[25] cpu_wdata[26]
+ cpu_wdata[27] cpu_wdata[28] cpu_wdata[29] cpu_wdata[2] cpu_wdata[30] cpu_wdata[31]
+ cpu_wdata[32] cpu_wdata[33] cpu_wdata[34] cpu_wdata[35] cpu_wdata[36] cpu_wdata[37]
+ cpu_wdata[38] cpu_wdata[39] cpu_wdata[3] cpu_wdata[40] cpu_wdata[41] cpu_wdata[42]
+ cpu_wdata[43] cpu_wdata[44] cpu_wdata[45] cpu_wdata[46] cpu_wdata[47] cpu_wdata[48]
+ cpu_wdata[49] cpu_wdata[4] cpu_wdata[50] cpu_wdata[51] cpu_wdata[52] cpu_wdata[53]
+ cpu_wdata[54] cpu_wdata[55] cpu_wdata[56] cpu_wdata[57] cpu_wdata[58] cpu_wdata[59]
+ cpu_wdata[5] cpu_wdata[60] cpu_wdata[61] cpu_wdata[62] cpu_wdata[63] cpu_wdata[6]
+ cpu_wdata[7] cpu_wdata[8] cpu_wdata[9] cpu_write mem_addr[0] mem_addr[10] mem_addr[11]
+ mem_addr[12] mem_addr[13] mem_addr[14] mem_addr[15] mem_addr[16] mem_addr[17] mem_addr[18]
+ mem_addr[19] mem_addr[1] mem_addr[20] mem_addr[21] mem_addr[22] mem_addr[23] mem_addr[24]
+ mem_addr[25] mem_addr[26] mem_addr[27] mem_addr[28] mem_addr[29] mem_addr[2] mem_addr[30]
+ mem_addr[31] mem_addr[3] mem_addr[4] mem_addr[5] mem_addr[6] mem_addr[7] mem_addr[8]
+ mem_addr[9] mem_rdata[0] mem_rdata[10] mem_rdata[11] mem_rdata[12] mem_rdata[13]
+ mem_rdata[14] mem_rdata[15] mem_rdata[16] mem_rdata[17] mem_rdata[18] mem_rdata[19]
+ mem_rdata[1] mem_rdata[20] mem_rdata[21] mem_rdata[22] mem_rdata[23] mem_rdata[24]
+ mem_rdata[25] mem_rdata[26] mem_rdata[27] mem_rdata[28] mem_rdata[29] mem_rdata[2]
+ mem_rdata[30] mem_rdata[31] mem_rdata[32] mem_rdata[33] mem_rdata[34] mem_rdata[35]
+ mem_rdata[36] mem_rdata[37] mem_rdata[38] mem_rdata[39] mem_rdata[3] mem_rdata[40]
+ mem_rdata[41] mem_rdata[42] mem_rdata[43] mem_rdata[44] mem_rdata[45] mem_rdata[46]
+ mem_rdata[47] mem_rdata[48] mem_rdata[49] mem_rdata[4] mem_rdata[50] mem_rdata[51]
+ mem_rdata[52] mem_rdata[53] mem_rdata[54] mem_rdata[55] mem_rdata[56] mem_rdata[57]
+ mem_rdata[58] mem_rdata[59] mem_rdata[5] mem_rdata[60] mem_rdata[61] mem_rdata[62]
+ mem_rdata[63] mem_rdata[6] mem_rdata[7] mem_rdata[8] mem_rdata[9] mem_read mem_ready
+ mem_wdata[0] mem_wdata[10] mem_wdata[11] mem_wdata[12] mem_wdata[13] mem_wdata[14]
+ mem_wdata[15] mem_wdata[16] mem_wdata[17] mem_wdata[18] mem_wdata[19] mem_wdata[1]
+ mem_wdata[20] mem_wdata[21] mem_wdata[22] mem_wdata[23] mem_wdata[24] mem_wdata[25]
+ mem_wdata[26] mem_wdata[27] mem_wdata[28] mem_wdata[29] mem_wdata[2] mem_wdata[30]
+ mem_wdata[31] mem_wdata[32] mem_wdata[33] mem_wdata[34] mem_wdata[35] mem_wdata[36]
+ mem_wdata[37] mem_wdata[38] mem_wdata[39] mem_wdata[3] mem_wdata[40] mem_wdata[41]
+ mem_wdata[42] mem_wdata[43] mem_wdata[44] mem_wdata[45] mem_wdata[46] mem_wdata[47]
+ mem_wdata[48] mem_wdata[49] mem_wdata[4] mem_wdata[50] mem_wdata[51] mem_wdata[52]
+ mem_wdata[53] mem_wdata[54] mem_wdata[55] mem_wdata[56] mem_wdata[57] mem_wdata[58]
+ mem_wdata[59] mem_wdata[5] mem_wdata[60] mem_wdata[61] mem_wdata[62] mem_wdata[63]
+ mem_wdata[6] mem_wdata[7] mem_wdata[8] mem_wdata[9] mem_write reset
XFILLER_100_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05903_ data_array.rdata0\[24\] net1666 net1147 VGND VGND VPWR VPWR _03396_ sky130_fd_sc_hd__o21a_1
X_06883_ data_array.data0\[0\]\[13\] net1363 net1269 data_array.data0\[3\]\[13\] _04174_
+ VGND VGND VPWR VPWR _04175_ sky130_fd_sc_hd__a221o_1
X_09671_ net704 net3522 net614 VGND VGND VPWR VPWR _01423_ sky130_fd_sc_hd__mux2_1
X_05834_ data_array.rdata0\[1\] net846 net1142 VGND VGND VPWR VPWR _03350_ sky130_fd_sc_hd__o21a_1
X_08622_ net734 net4316 net517 VGND VGND VPWR VPWR _00381_ sky130_fd_sc_hd__mux2_1
X_08553_ net742 net4423 net584 VGND VGND VPWR VPWR _00321_ sky130_fd_sc_hd__mux2_1
X_05765_ net4 fsm.tag_out1\[5\] VGND VGND VPWR VPWR _03282_ sky130_fd_sc_hd__xor2_2
XFILLER_51_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07504_ net1622 _04733_ _04737_ net1196 VGND VGND VPWR VPWR _04740_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_59_Left_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08484_ net824 net813 net855 _05558_ VGND VGND VPWR VPWR _05560_ sky130_fd_sc_hd__or4_1
XFILLER_22_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05696_ _03159_ _03212_ _03192_ _03177_ VGND VGND VPWR VPWR _03213_ sky130_fd_sc_hd__or4_4
XFILLER_161_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07435_ data_array.data0\[8\]\[63\] net1357 net1263 data_array.data0\[11\]\[63\]
+ _04676_ VGND VGND VPWR VPWR _04677_ sky130_fd_sc_hd__a221o_1
XFILLER_167_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07366_ data_array.data0\[1\]\[57\] net1538 net1442 data_array.data0\[2\]\[57\] VGND
+ VGND VPWR VPWR _04614_ sky130_fd_sc_hd__a22o_1
XFILLER_148_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09105_ net866 net3123 net413 VGND VGND VPWR VPWR _00859_ sky130_fd_sc_hd__mux2_1
X_06317_ net1229 _03655_ _03659_ net1181 VGND VGND VPWR VPWR _03661_ sky130_fd_sc_hd__a22o_1
XFILLER_149_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07297_ _04550_ _04551_ VGND VGND VPWR VPWR _00045_ sky130_fd_sc_hd__or2_1
XFILLER_136_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09036_ net2538 net881 net421 VGND VGND VPWR VPWR _00791_ sky130_fd_sc_hd__mux2_1
XFILLER_164_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06248_ tag_array.tag0\[1\]\[5\] net1607 net1511 tag_array.tag0\[2\]\[5\] VGND VGND
+ VPWR VPWR _03598_ sky130_fd_sc_hd__a22o_1
Xhold340 data_array.data0\[0\]\[41\] VGND VGND VPWR VPWR net1991 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_68_Left_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06179_ tag_array.valid1\[0\] net1366 net1272 tag_array.valid1\[3\] _03534_ VGND
+ VGND VPWR VPWR _03535_ sky130_fd_sc_hd__a221o_1
Xhold351 data_array.data1\[4\]\[2\] VGND VGND VPWR VPWR net2002 sky130_fd_sc_hd__dlygate4sd3_1
Xhold362 data_array.data1\[4\]\[9\] VGND VGND VPWR VPWR net2013 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold373 data_array.data0\[4\]\[48\] VGND VGND VPWR VPWR net2024 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold384 data_array.data1\[1\]\[11\] VGND VGND VPWR VPWR net2035 sky130_fd_sc_hd__dlygate4sd3_1
Xhold395 data_array.data0\[1\]\[63\] VGND VGND VPWR VPWR net2046 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout820 _05356_ VGND VGND VPWR VPWR net820 sky130_fd_sc_hd__buf_1
XFILLER_89_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout831 net835 VGND VGND VPWR VPWR net831 sky130_fd_sc_hd__buf_6
Xfanout842 net843 VGND VGND VPWR VPWR net842 sky130_fd_sc_hd__buf_6
X_09938_ net1076 net2883 net371 VGND VGND VPWR VPWR _01687_ sky130_fd_sc_hd__mux2_1
Xfanout853 _03213_ VGND VGND VPWR VPWR net853 sky130_fd_sc_hd__buf_12
Xfanout864 _05542_ VGND VGND VPWR VPWR net864 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_142_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout875 _05538_ VGND VGND VPWR VPWR net875 sky130_fd_sc_hd__clkbuf_2
XFILLER_133_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout886 _05532_ VGND VGND VPWR VPWR net886 sky130_fd_sc_hd__clkbuf_2
Xfanout897 _05526_ VGND VGND VPWR VPWR net897 sky130_fd_sc_hd__buf_1
X_09869_ net993 net4267 net383 VGND VGND VPWR VPWR _01619_ sky130_fd_sc_hd__mux2_1
Xhold1040 data_array.data1\[9\]\[7\] VGND VGND VPWR VPWR net2691 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1051 tag_array.tag0\[3\]\[24\] VGND VGND VPWR VPWR net2702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1062 tag_array.tag1\[10\]\[11\] VGND VGND VPWR VPWR net2713 sky130_fd_sc_hd__dlygate4sd3_1
X_11900_ clknet_leaf_89_clk _00708_ VGND VGND VPWR VPWR data_array.data0\[5\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1073 tag_array.tag1\[5\]\[16\] VGND VGND VPWR VPWR net2724 sky130_fd_sc_hd__dlygate4sd3_1
X_12880_ clknet_leaf_72_clk _01574_ VGND VGND VPWR VPWR data_array.data0\[12\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_172_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1084 data_array.data1\[0\]\[40\] VGND VGND VPWR VPWR net2735 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1095 tag_array.tag1\[10\]\[24\] VGND VGND VPWR VPWR net2746 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_77_Left_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11831_ clknet_leaf_90_clk _00639_ VGND VGND VPWR VPWR data_array.data0\[7\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_984 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11762_ clknet_leaf_31_clk _00570_ VGND VGND VPWR VPWR data_array.data0\[8\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13501_ clknet_leaf_29_clk _02130_ VGND VGND VPWR VPWR tag_array.dirty1\[0\] sky130_fd_sc_hd__dfxtp_1
X_10713_ net1813 net865 net482 VGND VGND VPWR VPWR _02458_ sky130_fd_sc_hd__mux2_1
X_14481_ clknet_leaf_161_clk _03104_ VGND VGND VPWR VPWR tag_array.dirty0\[15\] sky130_fd_sc_hd__dfxtp_1
X_11693_ clknet_leaf_127_clk _00501_ VGND VGND VPWR VPWR tag_array.tag1\[15\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13432_ clknet_leaf_209_clk _02062_ VGND VGND VPWR VPWR data_array.data1\[8\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
X_10644_ net2277 net886 net467 VGND VGND VPWR VPWR _02389_ sky130_fd_sc_hd__mux2_1
X_10575_ net907 net4442 net453 VGND VGND VPWR VPWR _02320_ sky130_fd_sc_hd__mux2_1
X_13363_ clknet_leaf_144_clk _01993_ VGND VGND VPWR VPWR tag_array.tag0\[2\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_127_536 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_86_Left_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12314_ clknet_leaf_102_clk _01072_ VGND VGND VPWR VPWR tag_array.tag1\[12\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13294_ clknet_leaf_47_clk _01924_ VGND VGND VPWR VPWR data_array.data0\[10\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_114_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12245_ clknet_leaf_31_clk _01003_ VGND VGND VPWR VPWR tag_array.tag1\[14\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_131_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12176_ clknet_leaf_145_clk _00984_ VGND VGND VPWR VPWR tag_array.tag0\[14\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_131_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11127_ net1010 net3129 net541 VGND VGND VPWR VPWR _02870_ sky130_fd_sc_hd__mux2_1
XFILLER_122_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11058_ net1841 net1028 net335 VGND VGND VPWR VPWR _02801_ sky130_fd_sc_hd__mux2_1
XFILLER_95_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10009_ net1050 net2886 net562 VGND VGND VPWR VPWR _01758_ sky130_fd_sc_hd__mux2_1
XFILLER_37_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_95_Left_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_177_3753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_177_3764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07220_ _04480_ _04481_ VGND VGND VPWR VPWR _00037_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_15_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07151_ data_array.data0\[4\]\[37\] net1355 net1261 data_array.data0\[7\]\[37\] _04418_
+ VGND VGND VPWR VPWR _04419_ sky130_fd_sc_hd__a221o_1
XFILLER_157_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06102_ data_array.rdata0\[17\] net1134 net1113 data_array.rdata1\[17\] VGND VGND
+ VPWR VPWR net271 sky130_fd_sc_hd__a22o_1
X_07082_ data_array.data0\[9\]\[31\] net1577 net1481 data_array.data0\[10\]\[31\]
+ VGND VGND VPWR VPWR _04356_ sky130_fd_sc_hd__a22o_1
XFILLER_172_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06033_ net1162 net1141 net1119 net28 VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__o31a_1
XFILLER_113_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07984_ data_array.data1\[9\]\[49\] net1572 net1476 data_array.data1\[10\]\[49\]
+ VGND VGND VPWR VPWR _05176_ sky130_fd_sc_hd__a22o_1
XFILLER_86_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09723_ net696 net3937 net611 VGND VGND VPWR VPWR _01475_ sky130_fd_sc_hd__mux2_1
XFILLER_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06935_ data_array.data0\[9\]\[18\] net1567 net1471 data_array.data0\[10\]\[18\]
+ VGND VGND VPWR VPWR _04222_ sky130_fd_sc_hd__a22o_1
XFILLER_101_469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09654_ net770 net4512 net614 VGND VGND VPWR VPWR _01406_ sky130_fd_sc_hd__mux2_1
X_06866_ net1628 _04153_ _04157_ net1202 VGND VGND VPWR VPWR _04160_ sky130_fd_sc_hd__a22o_1
X_08605_ net703 net3143 net528 VGND VGND VPWR VPWR _00364_ sky130_fd_sc_hd__mux2_1
XFILLER_82_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05817_ _03239_ _03277_ _03289_ VGND VGND VPWR VPWR _03334_ sky130_fd_sc_hd__or3_1
XFILLER_103_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09585_ net1010 net2765 net394 VGND VGND VPWR VPWR _01337_ sky130_fd_sc_hd__mux2_1
X_06797_ data_array.data0\[12\]\[5\] net1360 net1266 data_array.data0\[15\]\[5\] _04096_
+ VGND VGND VPWR VPWR _04097_ sky130_fd_sc_hd__a221o_1
XFILLER_63_17 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08536_ net814 _05561_ net1697 VGND VGND VPWR VPWR _00307_ sky130_fd_sc_hd__a21o_1
X_05748_ net9 fsm.tag_out1\[10\] VGND VGND VPWR VPWR _03265_ sky130_fd_sc_hd__and2b_1
XFILLER_179_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08467_ net814 _05547_ VGND VGND VPWR VPWR _05548_ sky130_fd_sc_hd__nand2_2
X_05679_ fsm.tag_out0\[6\] net5 VGND VGND VPWR VPWR _03196_ sky130_fd_sc_hd__and2b_1
X_07418_ _04660_ _04661_ VGND VGND VPWR VPWR _00057_ sky130_fd_sc_hd__or2_1
X_08398_ net1123 _05501_ VGND VGND VPWR VPWR _05502_ sky130_fd_sc_hd__and2_1
XFILLER_10_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_98_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07349_ data_array.data0\[4\]\[55\] net1343 net1249 data_array.data0\[7\]\[55\] _04598_
+ VGND VGND VPWR VPWR _04599_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_59_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10360_ net758 net2438 net540 VGND VGND VPWR VPWR _02107_ sky130_fd_sc_hd__mux2_1
XFILLER_124_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09019_ net3724 net948 net424 VGND VGND VPWR VPWR _00774_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_76_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10291_ net2176 net997 net635 VGND VGND VPWR VPWR _02038_ sky130_fd_sc_hd__mux2_1
X_12030_ clknet_leaf_109_clk _00838_ VGND VGND VPWR VPWR data_array.data0\[6\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_151_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold170 data_array.data1\[2\]\[53\] VGND VGND VPWR VPWR net1821 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 data_array.data1\[4\]\[58\] VGND VGND VPWR VPWR net1832 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 data_array.data1\[4\]\[26\] VGND VGND VPWR VPWR net1843 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout1604 net1606 VGND VGND VPWR VPWR net1604 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_72_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1615 net1617 VGND VGND VPWR VPWR net1615 sky130_fd_sc_hd__clkbuf_2
Xfanout1626 net1627 VGND VGND VPWR VPWR net1626 sky130_fd_sc_hd__clkbuf_4
XFILLER_137_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1637 _03506_ VGND VGND VPWR VPWR net1637 sky130_fd_sc_hd__buf_4
Xfanout650 net651 VGND VGND VPWR VPWR net650 sky130_fd_sc_hd__buf_4
Xfanout1648 net98 VGND VGND VPWR VPWR net1648 sky130_fd_sc_hd__buf_4
Xfanout661 net666 VGND VGND VPWR VPWR net661 sky130_fd_sc_hd__buf_4
Xfanout672 _05549_ VGND VGND VPWR VPWR net672 sky130_fd_sc_hd__buf_4
XFILLER_144_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout683 net684 VGND VGND VPWR VPWR net683 sky130_fd_sc_hd__buf_4
X_13981_ clknet_leaf_229_clk _02610_ VGND VGND VPWR VPWR data_array.data1\[5\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout694 net697 VGND VGND VPWR VPWR net694 sky130_fd_sc_hd__clkbuf_2
XFILLER_93_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_670 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12932_ clknet_leaf_85_clk _01626_ VGND VGND VPWR VPWR data_array.data0\[13\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12863_ clknet_leaf_34_clk _01557_ VGND VGND VPWR VPWR data_array.data0\[12\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11814_ clknet_leaf_223_clk _00622_ VGND VGND VPWR VPWR data_array.data0\[7\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_57_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12794_ clknet_leaf_167_clk _01488_ VGND VGND VPWR VPWR tag_array.tag1\[10\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_159_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11745_ clknet_leaf_45_clk _00553_ VGND VGND VPWR VPWR data_array.data0\[8\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_155_3336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14464_ clknet_leaf_73_clk _03087_ VGND VGND VPWR VPWR data_array.data1\[7\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_12_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11676_ clknet_leaf_129_clk _00484_ VGND VGND VPWR VPWR tag_array.tag1\[1\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_12_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13415_ clknet_leaf_259_clk _02045_ VGND VGND VPWR VPWR data_array.data1\[8\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
X_10627_ net2385 net952 net467 VGND VGND VPWR VPWR _02372_ sky130_fd_sc_hd__mux2_1
X_14395_ clknet_leaf_27_clk _03018_ VGND VGND VPWR VPWR data_array.data1\[10\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_133_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13346_ clknet_leaf_13_clk _01976_ VGND VGND VPWR VPWR data_array.data0\[10\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_127_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10558_ net975 net2427 net455 VGND VGND VPWR VPWR _02303_ sky130_fd_sc_hd__mux2_1
XFILLER_143_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13277_ clknet_leaf_241_clk _01907_ VGND VGND VPWR VPWR data_array.data0\[11\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_170_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10489_ net989 net3248 net349 VGND VGND VPWR VPWR _02234_ sky130_fd_sc_hd__mux2_1
X_12228_ clknet_leaf_148_clk _00157_ VGND VGND VPWR VPWR fsm.tag_out1\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_130_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12159_ clknet_leaf_157_clk _00967_ VGND VGND VPWR VPWR tag_array.tag0\[13\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_151_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1809 tag_array.tag1\[14\]\[15\] VGND VGND VPWR VPWR net3460 sky130_fd_sc_hd__dlygate4sd3_1
X_06720_ tag_array.tag1\[12\]\[23\] net1419 net1325 tag_array.tag1\[15\]\[23\] _04026_
+ VGND VGND VPWR VPWR _04027_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_179_3804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06651_ tag_array.tag1\[5\]\[17\] net1607 net1511 tag_array.tag1\[6\]\[17\] VGND
+ VGND VPWR VPWR _03964_ sky130_fd_sc_hd__a22o_1
XFILLER_25_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09370_ net920 net4472 net406 VGND VGND VPWR VPWR _01123_ sky130_fd_sc_hd__mux2_1
X_06582_ _03900_ _03901_ VGND VGND VPWR VPWR _00157_ sky130_fd_sc_hd__or2_2
X_08321_ net1753 net1048 net691 VGND VGND VPWR VPWR _00236_ sky130_fd_sc_hd__mux2_1
XFILLER_71_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08252_ fsm.tag_out1\[19\] net817 net809 fsm.tag_out0\[19\] _05402_ VGND VGND VPWR
+ VPWR _05403_ sky130_fd_sc_hd__a221o_1
XFILLER_177_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07203_ data_array.data0\[13\]\[42\] net1586 net1490 data_array.data0\[14\]\[42\]
+ VGND VGND VPWR VPWR _04466_ sky130_fd_sc_hd__a22o_1
X_08183_ _03511_ _03519_ net821 VGND VGND VPWR VPWR _05354_ sky130_fd_sc_hd__or3_1
Xclkbuf_4_12_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_12_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_31_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07134_ data_array.data0\[8\]\[36\] net1413 net1319 data_array.data0\[11\]\[36\]
+ _04402_ VGND VGND VPWR VPWR _04403_ sky130_fd_sc_hd__a221o_1
XFILLER_174_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07065_ net1225 _04335_ _04339_ net1178 VGND VGND VPWR VPWR _04341_ sky130_fd_sc_hd__a22o_1
XFILLER_134_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput220 net220 VGND VGND VPWR VPWR cpu_rdata[5] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_93_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput231 net231 VGND VGND VPWR VPWR mem_addr[10] sky130_fd_sc_hd__buf_2
X_06016_ net156 net1152 _03470_ _03471_ VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__a22o_1
Xoutput242 net242 VGND VGND VPWR VPWR mem_addr[20] sky130_fd_sc_hd__buf_2
Xoutput253 net253 VGND VGND VPWR VPWR mem_addr[30] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput264 net264 VGND VGND VPWR VPWR mem_wdata[10] sky130_fd_sc_hd__buf_2
XFILLER_114_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput275 net275 VGND VGND VPWR VPWR mem_wdata[20] sky130_fd_sc_hd__buf_2
Xoutput286 net286 VGND VGND VPWR VPWR mem_wdata[30] sky130_fd_sc_hd__buf_2
Xoutput297 net297 VGND VGND VPWR VPWR mem_wdata[40] sky130_fd_sc_hd__buf_2
X_07967_ net1180 _05155_ _05159_ net1228 VGND VGND VPWR VPWR _05161_ sky130_fd_sc_hd__a22o_1
X_09706_ net763 net4604 net611 VGND VGND VPWR VPWR _01458_ sky130_fd_sc_hd__mux2_1
X_06918_ data_array.data0\[12\]\[16\] net1356 net1262 data_array.data0\[15\]\[16\]
+ _04206_ VGND VGND VPWR VPWR _04207_ sky130_fd_sc_hd__a221o_1
X_07898_ data_array.data1\[1\]\[41\] net1525 net1429 data_array.data1\[2\]\[41\] VGND
+ VGND VPWR VPWR _05098_ sky130_fd_sc_hd__a22o_1
XFILLER_55_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09637_ net738 net2649 net617 VGND VGND VPWR VPWR _01389_ sky130_fd_sc_hd__mux2_1
XFILLER_16_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06849_ data_array.data0\[5\]\[10\] net1601 net1505 data_array.data0\[6\]\[10\] VGND
+ VGND VPWR VPWR _04144_ sky130_fd_sc_hd__a22o_1
XFILLER_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09568_ net1077 net3020 net395 VGND VGND VPWR VPWR _01320_ sky130_fd_sc_hd__mux2_1
XFILLER_70_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08519_ _03516_ _03519_ net823 VGND VGND VPWR VPWR _05584_ sky130_fd_sc_hd__or3_1
XFILLER_169_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09499_ net732 net4076 net625 VGND VGND VPWR VPWR _01252_ sky130_fd_sc_hd__mux2_1
X_11530_ clknet_leaf_175_clk _00338_ VGND VGND VPWR VPWR tag_array.valid1\[2\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_137_Right_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_478 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11461_ clknet_leaf_241_clk _00271_ VGND VGND VPWR VPWR data_array.data0\[0\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13200_ clknet_leaf_214_clk _00094_ VGND VGND VPWR VPWR data_array.rdata1\[37\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_150_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10412_ net1774 net1004 net662 VGND VGND VPWR VPWR _02158_ sky130_fd_sc_hd__mux2_1
XFILLER_136_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_150_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11392_ clknet_leaf_189_clk _00202_ VGND VGND VPWR VPWR tag_array.tag1\[7\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_14180_ clknet_leaf_26_clk _02809_ VGND VGND VPWR VPWR data_array.data0\[2\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13131_ clknet_leaf_180_clk _01825_ VGND VGND VPWR VPWR tag_array.tag0\[3\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_109_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10343_ net726 net3629 net593 VGND VGND VPWR VPWR _02090_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_111_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13062_ clknet_leaf_200_clk _01756_ VGND VGND VPWR VPWR data_array.data1\[13\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_10274_ net1796 net1067 net644 VGND VGND VPWR VPWR _02021_ sky130_fd_sc_hd__mux2_1
XFILLER_151_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12013_ clknet_leaf_175_clk _00821_ VGND VGND VPWR VPWR data_array.data0\[6\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_79_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1401 net1403 VGND VGND VPWR VPWR net1401 sky130_fd_sc_hd__clkbuf_4
Xfanout1412 net1413 VGND VGND VPWR VPWR net1412 sky130_fd_sc_hd__clkbuf_4
Xfanout1423 net1425 VGND VGND VPWR VPWR net1423 sky130_fd_sc_hd__clkbuf_4
Xfanout1434 net1447 VGND VGND VPWR VPWR net1434 sky130_fd_sc_hd__clkbuf_2
Xfanout1445 net1446 VGND VGND VPWR VPWR net1445 sky130_fd_sc_hd__clkbuf_4
XFILLER_78_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1456 net1458 VGND VGND VPWR VPWR net1456 sky130_fd_sc_hd__clkbuf_4
Xfanout1467 net1470 VGND VGND VPWR VPWR net1467 sky130_fd_sc_hd__clkbuf_2
XFILLER_171_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout480 net489 VGND VGND VPWR VPWR net480 sky130_fd_sc_hd__buf_4
Xfanout1478 net1480 VGND VGND VPWR VPWR net1478 sky130_fd_sc_hd__clkbuf_4
Xfanout491 net495 VGND VGND VPWR VPWR net491 sky130_fd_sc_hd__buf_2
XFILLER_87_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1489 net1491 VGND VGND VPWR VPWR net1489 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13964_ clknet_leaf_68_clk _02593_ VGND VGND VPWR VPWR data_array.data1\[5\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_109_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12915_ clknet_leaf_60_clk _01609_ VGND VGND VPWR VPWR data_array.data0\[13\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13895_ clknet_leaf_193_clk _02524_ VGND VGND VPWR VPWR data_array.data1\[3\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_17_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12846_ clknet_leaf_51_clk _01540_ VGND VGND VPWR VPWR data_array.data0\[12\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_181_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12777_ clknet_leaf_169_clk _01471_ VGND VGND VPWR VPWR tag_array.tag0\[6\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_14_Left_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11728_ clknet_leaf_161_clk _00536_ VGND VGND VPWR VPWR tag_array.tag0\[9\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_147_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_104_Right_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14447_ clknet_leaf_37_clk _03070_ VGND VGND VPWR VPWR data_array.data1\[7\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_11659_ clknet_leaf_97_clk _00467_ VGND VGND VPWR VPWR tag_array.tag1\[1\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_156_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14378_ clknet_leaf_31_clk _03001_ VGND VGND VPWR VPWR data_array.data1\[10\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_155_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold906 data_array.data0\[4\]\[54\] VGND VGND VPWR VPWR net2557 sky130_fd_sc_hd__dlygate4sd3_1
Xhold917 tag_array.dirty1\[2\] VGND VGND VPWR VPWR net2568 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13329_ clknet_leaf_73_clk _01959_ VGND VGND VPWR VPWR data_array.data0\[10\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold928 tag_array.tag0\[3\]\[22\] VGND VGND VPWR VPWR net2579 sky130_fd_sc_hd__dlygate4sd3_1
Xhold939 data_array.data1\[14\]\[13\] VGND VGND VPWR VPWR net2590 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_50_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2307 data_array.data0\[10\]\[14\] VGND VGND VPWR VPWR net3958 sky130_fd_sc_hd__dlygate4sd3_1
X_08870_ net1026 net4164 net437 VGND VGND VPWR VPWR _00627_ sky130_fd_sc_hd__mux2_1
Xhold2318 data_array.data1\[9\]\[33\] VGND VGND VPWR VPWR net3969 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2329 tag_array.tag1\[7\]\[7\] VGND VGND VPWR VPWR net3980 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07821_ data_array.data1\[1\]\[34\] net1531 net1435 data_array.data1\[2\]\[34\] VGND
+ VGND VPWR VPWR _05028_ sky130_fd_sc_hd__a22o_1
Xhold1606 tag_array.tag0\[7\]\[19\] VGND VGND VPWR VPWR net3257 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1617 tag_array.tag0\[10\]\[14\] VGND VGND VPWR VPWR net3268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1628 data_array.data0\[11\]\[19\] VGND VGND VPWR VPWR net3279 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1639 data_array.data1\[2\]\[24\] VGND VGND VPWR VPWR net3290 sky130_fd_sc_hd__dlygate4sd3_1
X_07752_ data_array.data1\[4\]\[28\] net1349 net1255 data_array.data1\[7\]\[28\] _04964_
+ VGND VGND VPWR VPWR _04965_ sky130_fd_sc_hd__a221o_1
XFILLER_37_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06703_ _04010_ _04011_ VGND VGND VPWR VPWR _00169_ sky130_fd_sc_hd__or2_1
X_07683_ data_array.data1\[9\]\[22\] net1537 net1441 data_array.data1\[10\]\[22\]
+ VGND VGND VPWR VPWR _04902_ sky130_fd_sc_hd__a22o_1
XFILLER_53_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09422_ net979 net3969 net586 VGND VGND VPWR VPWR _01175_ sky130_fd_sc_hd__mux2_1
X_06634_ tag_array.tag1\[4\]\[15\] net1388 net1294 tag_array.tag1\[7\]\[15\] _03948_
+ VGND VGND VPWR VPWR _03949_ sky130_fd_sc_hd__a221o_1
XFILLER_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09353_ net988 net3903 net407 VGND VGND VPWR VPWR _01106_ sky130_fd_sc_hd__mux2_1
X_06565_ tag_array.tag1\[13\]\[9\] net1609 net1513 tag_array.tag1\[14\]\[9\] VGND
+ VGND VPWR VPWR _03886_ sky130_fd_sc_hd__a22o_1
XFILLER_178_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08304_ net100 net35 net1648 VGND VGND VPWR VPWR _05439_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06496_ tag_array.tag1\[8\]\[3\] net1372 net1278 tag_array.tag1\[11\]\[3\] _03822_
+ VGND VGND VPWR VPWR _03823_ sky130_fd_sc_hd__a221o_1
X_09284_ net742 net4140 net559 VGND VGND VPWR VPWR _01038_ sky130_fd_sc_hd__mux2_1
XFILLER_166_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08235_ net740 net2919 net805 VGND VGND VPWR VPWR _00209_ sky130_fd_sc_hd__mux2_1
XFILLER_166_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08166_ _05340_ _05341_ VGND VGND VPWR VPWR _00129_ sky130_fd_sc_hd__or2_1
XFILLER_118_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07117_ data_array.data0\[1\]\[34\] net1531 net1435 data_array.data0\[2\]\[34\] VGND
+ VGND VPWR VPWR _04388_ sky130_fd_sc_hd__a22o_1
X_08097_ data_array.data1\[4\]\[59\] net1379 net1285 data_array.data1\[7\]\[59\] _05278_
+ VGND VGND VPWR VPWR _05279_ sky130_fd_sc_hd__a221o_1
XFILLER_134_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07048_ data_array.data0\[4\]\[28\] net1350 net1256 data_array.data0\[7\]\[28\] _04324_
+ VGND VGND VPWR VPWR _04325_ sky130_fd_sc_hd__a221o_1
Xclkload90 clknet_leaf_62_clk VGND VGND VPWR VPWR clkload90/Y sky130_fd_sc_hd__bufinv_16
XFILLER_121_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2830 data_array.data0\[11\]\[14\] VGND VGND VPWR VPWR net4481 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2841 data_array.data0\[13\]\[50\] VGND VGND VPWR VPWR net4492 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2852 data_array.data1\[10\]\[0\] VGND VGND VPWR VPWR net4503 sky130_fd_sc_hd__dlygate4sd3_1
X_08999_ net2786 net1028 net424 VGND VGND VPWR VPWR _00754_ sky130_fd_sc_hd__mux2_1
XFILLER_85_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2863 data_array.data1\[15\]\[37\] VGND VGND VPWR VPWR net4514 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2874 data_array.data0\[15\]\[39\] VGND VGND VPWR VPWR net4525 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2885 data_array.data1\[11\]\[51\] VGND VGND VPWR VPWR net4536 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2896 data_array.data0\[3\]\[3\] VGND VGND VPWR VPWR net4547 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10961_ net898 net3403 net530 VGND VGND VPWR VPWR _02706_ sky130_fd_sc_hd__mux2_1
XFILLER_16_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_470 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12700_ clknet_leaf_182_clk _01394_ VGND VGND VPWR VPWR tag_array.tag0\[8\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_13680_ clknet_leaf_122_clk _02309_ VGND VGND VPWR VPWR data_array.data1\[15\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_55_194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10892_ net918 net3321 net520 VGND VGND VPWR VPWR _02637_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12631_ clknet_leaf_192_clk _01325_ VGND VGND VPWR VPWR data_array.data0\[15\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_43_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12562_ clknet_leaf_161_clk _01256_ VGND VGND VPWR VPWR tag_array.tag0\[11\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1018 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14301_ clknet_leaf_228_clk _02930_ VGND VGND VPWR VPWR data_array.data1\[11\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_11513_ clknet_leaf_167_clk _00321_ VGND VGND VPWR VPWR tag_array.tag1\[9\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12493_ clknet_leaf_27_clk _01187_ VGND VGND VPWR VPWR data_array.data1\[9\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
X_14232_ clknet_leaf_213_clk _02861_ VGND VGND VPWR VPWR data_array.data1\[12\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_11444_ clknet_leaf_89_clk _00254_ VGND VGND VPWR VPWR data_array.data0\[0\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14163_ clknet_leaf_43_clk _02792_ VGND VGND VPWR VPWR data_array.data0\[2\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_11375_ net819 net3583 _05584_ VGND VGND VPWR VPWR _03118_ sky130_fd_sc_hd__mux2_1
XFILLER_125_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13114_ clknet_leaf_166_clk _01808_ VGND VGND VPWR VPWR tag_array.tag0\[3\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_180_773 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10326_ net2560 net859 net637 VGND VGND VPWR VPWR _02073_ sky130_fd_sc_hd__mux2_1
X_14094_ clknet_leaf_1_clk _02723_ VGND VGND VPWR VPWR data_array.data0\[1\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_112_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_167_3571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ clknet_leaf_110_clk _01739_ VGND VGND VPWR VPWR data_array.data0\[3\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
X_10257_ net717 net2466 net596 VGND VGND VPWR VPWR _02004_ sky130_fd_sc_hd__mux2_1
Xfanout1220 net1223 VGND VGND VPWR VPWR net1220 sky130_fd_sc_hd__buf_2
XFILLER_39_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1231 net1233 VGND VGND VPWR VPWR net1231 sky130_fd_sc_hd__buf_4
XFILLER_182_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1242 net1245 VGND VGND VPWR VPWR net1242 sky130_fd_sc_hd__clkbuf_4
X_10188_ net1053 net3958 net358 VGND VGND VPWR VPWR _01935_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1253 net1254 VGND VGND VPWR VPWR net1253 sky130_fd_sc_hd__clkbuf_4
XFILLER_66_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1264 net1270 VGND VGND VPWR VPWR net1264 sky130_fd_sc_hd__clkbuf_2
XFILLER_78_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1275 net1276 VGND VGND VPWR VPWR net1275 sky130_fd_sc_hd__clkbuf_4
XFILLER_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1286 net1288 VGND VGND VPWR VPWR net1286 sky130_fd_sc_hd__clkbuf_2
XFILLER_93_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1297 net1298 VGND VGND VPWR VPWR net1297 sky130_fd_sc_hd__clkbuf_4
X_13947_ clknet_leaf_4_clk _02576_ VGND VGND VPWR VPWR data_array.data1\[4\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_868 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13878_ clknet_leaf_261_clk _02507_ VGND VGND VPWR VPWR data_array.data1\[3\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_22_Left_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12829_ clknet_leaf_196_clk _01523_ VGND VGND VPWR VPWR tag_array.tag1\[0\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06350_ net1173 _03685_ _03689_ net1222 VGND VGND VPWR VPWR _03691_ sky130_fd_sc_hd__a22o_1
XFILLER_91_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06281_ tag_array.tag0\[5\]\[8\] net1598 net1502 tag_array.tag0\[6\]\[8\] VGND VGND
+ VPWR VPWR _03628_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_150_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_150_clk
+ sky130_fd_sc_hd__clkbuf_8
X_08020_ data_array.data1\[0\]\[52\] net1354 net1260 data_array.data1\[3\]\[52\] _05208_
+ VGND VGND VPWR VPWR _05209_ sky130_fd_sc_hd__a221o_1
XFILLER_175_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold703 data_array.data0\[6\]\[47\] VGND VGND VPWR VPWR net2354 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_932 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold714 data_array.data1\[8\]\[8\] VGND VGND VPWR VPWR net2365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold725 data_array.data0\[1\]\[52\] VGND VGND VPWR VPWR net2376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold736 data_array.data1\[7\]\[13\] VGND VGND VPWR VPWR net2387 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_31_Left_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold747 data_array.data1\[2\]\[16\] VGND VGND VPWR VPWR net2398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold758 data_array.data0\[15\]\[10\] VGND VGND VPWR VPWR net2409 sky130_fd_sc_hd__dlygate4sd3_1
X_09971_ net945 net4283 net370 VGND VGND VPWR VPWR _01720_ sky130_fd_sc_hd__mux2_1
Xhold769 tag_array.dirty0\[13\] VGND VGND VPWR VPWR net2420 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_626 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08922_ net1076 net3226 net426 VGND VGND VPWR VPWR _00678_ sky130_fd_sc_hd__mux2_1
XFILLER_69_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2104 data_array.data0\[6\]\[54\] VGND VGND VPWR VPWR net3755 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2115 tag_array.tag0\[13\]\[5\] VGND VGND VPWR VPWR net3766 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2126 tag_array.tag1\[3\]\[1\] VGND VGND VPWR VPWR net3777 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2137 data_array.data0\[9\]\[15\] VGND VGND VPWR VPWR net3788 sky130_fd_sc_hd__dlygate4sd3_1
X_08853_ net1092 net3837 net439 VGND VGND VPWR VPWR _00610_ sky130_fd_sc_hd__mux2_1
Xhold2148 data_array.data1\[15\]\[61\] VGND VGND VPWR VPWR net3799 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1403 data_array.data1\[15\]\[45\] VGND VGND VPWR VPWR net3054 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1414 data_array.data1\[7\]\[5\] VGND VGND VPWR VPWR net3065 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2159 data_array.data1\[6\]\[11\] VGND VGND VPWR VPWR net3810 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1425 data_array.data1\[12\]\[57\] VGND VGND VPWR VPWR net3076 sky130_fd_sc_hd__dlygate4sd3_1
X_07804_ data_array.data1\[13\]\[33\] net1588 net1492 data_array.data1\[14\]\[33\]
+ VGND VGND VPWR VPWR _05012_ sky130_fd_sc_hd__a22o_1
Xhold1436 data_array.data0\[10\]\[10\] VGND VGND VPWR VPWR net3087 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1447 data_array.data0\[14\]\[54\] VGND VGND VPWR VPWR net3098 sky130_fd_sc_hd__dlygate4sd3_1
X_08784_ net3207 net1108 net445 VGND VGND VPWR VPWR _00542_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1458 data_array.data0\[15\]\[41\] VGND VGND VPWR VPWR net3109 sky130_fd_sc_hd__dlygate4sd3_1
X_05996_ data_array.rdata0\[55\] net853 net1146 VGND VGND VPWR VPWR _03458_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_88_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1469 data_array.data1\[13\]\[18\] VGND VGND VPWR VPWR net3120 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_0_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07735_ net1616 _04943_ _04947_ net1190 VGND VGND VPWR VPWR _04950_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_49_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Left_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07666_ data_array.data1\[8\]\[20\] net1419 net1325 data_array.data1\[11\]\[20\]
+ _04886_ VGND VGND VPWR VPWR _04887_ sky130_fd_sc_hd__a221o_1
XFILLER_41_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09405_ net1044 net3754 net582 VGND VGND VPWR VPWR _01158_ sky130_fd_sc_hd__mux2_1
XFILLER_164_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06617_ tag_array.tag1\[8\]\[14\] net1368 net1274 tag_array.tag1\[11\]\[14\] _03932_
+ VGND VGND VPWR VPWR _03933_ sky130_fd_sc_hd__a221o_1
XFILLER_111_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07597_ data_array.data1\[5\]\[14\] net1570 net1474 data_array.data1\[6\]\[14\] VGND
+ VGND VPWR VPWR _04824_ sky130_fd_sc_hd__a22o_1
X_09336_ net1059 net3530 net404 VGND VGND VPWR VPWR _01089_ sky130_fd_sc_hd__mux2_1
X_06548_ net1185 _03865_ _03869_ net1233 VGND VGND VPWR VPWR _03871_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_62_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09267_ net710 net3034 net569 VGND VGND VPWR VPWR _01021_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_141_clk clknet_5_31__leaf_clk VGND VGND VPWR VPWR clknet_leaf_141_clk
+ sky130_fd_sc_hd__clkbuf_8
X_06479_ tag_array.tag1\[1\]\[1\] net1575 net1479 tag_array.tag1\[2\]\[1\] VGND VGND
+ VPWR VPWR _03808_ sky130_fd_sc_hd__a22o_1
X_08218_ net1650 net1162 net7 VGND VGND VPWR VPWR _05380_ sky130_fd_sc_hd__and3_1
XFILLER_154_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09198_ net790 net3596 net630 VGND VGND VPWR VPWR _00952_ sky130_fd_sc_hd__mux2_1
XFILLER_14_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08149_ tag_array.dirty1\[9\] net1574 net1478 tag_array.dirty1\[10\] VGND VGND VPWR
+ VPWR _05326_ sky130_fd_sc_hd__a22o_1
XFILLER_119_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11160_ net879 net3196 net545 VGND VGND VPWR VPWR _02903_ sky130_fd_sc_hd__mux2_1
Xclkload190 clknet_leaf_99_clk VGND VGND VPWR VPWR clkload190/Y sky130_fd_sc_hd__bufinv_16
X_10111_ net1103 net2900 net364 VGND VGND VPWR VPWR _01859_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11091_ net2085 net896 net328 VGND VGND VPWR VPWR _02834_ sky130_fd_sc_hd__mux2_1
XFILLER_96_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10042_ net918 net2977 net562 VGND VGND VPWR VPWR _01791_ sky130_fd_sc_hd__mux2_1
XFILLER_1_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_145_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2660 tag_array.tag1\[3\]\[15\] VGND VGND VPWR VPWR net4311 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 tag_array.valid0\[6\] VGND VGND VPWR VPWR net1703 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2671 data_array.data1\[3\]\[24\] VGND VGND VPWR VPWR net4322 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_69_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold63 tag_array.valid0\[7\] VGND VGND VPWR VPWR net1714 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold74 data_array.data1\[1\]\[15\] VGND VGND VPWR VPWR net1725 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2682 tag_array.tag0\[4\]\[4\] VGND VGND VPWR VPWR net4333 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 data_array.data1\[1\]\[60\] VGND VGND VPWR VPWR net1736 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2693 tag_array.tag0\[5\]\[17\] VGND VGND VPWR VPWR net4344 sky130_fd_sc_hd__dlygate4sd3_1
X_13801_ clknet_leaf_73_clk _02430_ VGND VGND VPWR VPWR data_array.data1\[2\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold96 tag_array.tag1\[2\]\[22\] VGND VGND VPWR VPWR net1747 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1970 tag_array.tag0\[14\]\[19\] VGND VGND VPWR VPWR net3621 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1981 tag_array.tag0\[2\]\[6\] VGND VGND VPWR VPWR net3632 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1992 data_array.data1\[14\]\[27\] VGND VGND VPWR VPWR net3643 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_63_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11993_ clknet_leaf_49_clk _00801_ VGND VGND VPWR VPWR data_array.data0\[6\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13732_ clknet_leaf_234_clk _02361_ VGND VGND VPWR VPWR data_array.data1\[1\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_10944_ net966 net2799 net535 VGND VGND VPWR VPWR _02689_ sky130_fd_sc_hd__mux2_1
XFILLER_16_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13663_ clknet_leaf_204_clk _02292_ VGND VGND VPWR VPWR data_array.data1\[15\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10875_ net984 net3221 net519 VGND VGND VPWR VPWR _02620_ sky130_fd_sc_hd__mux2_1
X_12614_ clknet_leaf_156_clk _01308_ VGND VGND VPWR VPWR tag_array.tag0\[0\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_169_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13594_ clknet_leaf_60_clk _02223_ VGND VGND VPWR VPWR data_array.data0\[9\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_12545_ clknet_leaf_170_clk _01239_ VGND VGND VPWR VPWR tag_array.tag0\[11\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_132_clk clknet_5_30__leaf_clk VGND VGND VPWR VPWR clknet_leaf_132_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_40_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12476_ clknet_leaf_31_clk _01170_ VGND VGND VPWR VPWR data_array.data1\[9\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_169_3600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14215_ clknet_leaf_224_clk _02844_ VGND VGND VPWR VPWR data_array.data0\[2\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_169_3611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11427_ clknet_leaf_222_clk _00237_ VGND VGND VPWR VPWR data_array.data0\[0\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_5 _00107_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14146_ clknet_leaf_208_clk _02775_ VGND VGND VPWR VPWR data_array.data0\[1\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
X_11358_ net862 net3663 net804 VGND VGND VPWR VPWR _03101_ sky130_fd_sc_hd__mux2_1
XFILLER_113_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10309_ net1967 net925 net633 VGND VGND VPWR VPWR _02056_ sky130_fd_sc_hd__mux2_1
X_14077_ clknet_leaf_3_clk _02706_ VGND VGND VPWR VPWR data_array.data1\[6\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11289_ net874 net4165 net680 VGND VGND VPWR VPWR _03032_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_182_3855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13028_ clknet_leaf_49_clk _01722_ VGND VGND VPWR VPWR data_array.data0\[3\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_199_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_199_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_67_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1050 net1051 VGND VGND VPWR VPWR net1050 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1061 _05444_ VGND VGND VPWR VPWR net1061 sky130_fd_sc_hd__dlymetal6s2s_1
X_05850_ data_array.rdata1\[6\] net828 net837 VGND VGND VPWR VPWR _03361_ sky130_fd_sc_hd__a21o_1
Xfanout1072 _05438_ VGND VGND VPWR VPWR net1072 sky130_fd_sc_hd__clkbuf_2
Xfanout1083 _05434_ VGND VGND VPWR VPWR net1083 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1094 _05428_ VGND VGND VPWR VPWR net1094 sky130_fd_sc_hd__clkbuf_2
XFILLER_66_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05781_ fsm.tag_out1\[11\] net10 VGND VGND VPWR VPWR _03298_ sky130_fd_sc_hd__and2b_1
X_07520_ data_array.data1\[1\]\[7\] net1589 net1493 data_array.data1\[2\]\[7\] VGND
+ VGND VPWR VPWR _04754_ sky130_fd_sc_hd__a22o_1
XFILLER_179_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07451_ _04690_ _04691_ VGND VGND VPWR VPWR _00064_ sky130_fd_sc_hd__or2_1
X_06402_ tag_array.tag0\[5\]\[19\] net1596 net1500 tag_array.tag0\[6\]\[19\] VGND
+ VGND VPWR VPWR _03738_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_44_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07382_ data_array.data0\[0\]\[58\] net1355 net1261 data_array.data0\[3\]\[58\] _04628_
+ VGND VGND VPWR VPWR _04629_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_44_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_106_Left_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09121_ net1057 net2590 net570 VGND VGND VPWR VPWR _00875_ sky130_fd_sc_hd__mux2_1
X_06333_ tag_array.tag0\[0\]\[13\] net1417 net1323 tag_array.tag0\[3\]\[13\] _03674_
+ VGND VGND VPWR VPWR _03675_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_123_clk clknet_5_27__leaf_clk VGND VGND VPWR VPWR clknet_leaf_123_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_175_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09052_ net1076 net3024 net410 VGND VGND VPWR VPWR _00806_ sky130_fd_sc_hd__mux2_1
X_06264_ tag_array.tag0\[9\]\[7\] net1598 net1502 tag_array.tag0\[10\]\[7\] VGND VGND
+ VPWR VPWR _03612_ sky130_fd_sc_hd__a22o_1
XFILLER_148_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08003_ data_array.data1\[12\]\[51\] net1333 net1239 data_array.data1\[15\]\[51\]
+ _05192_ VGND VGND VPWR VPWR _05193_ sky130_fd_sc_hd__a221o_1
XFILLER_163_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold500 data_array.data0\[0\]\[53\] VGND VGND VPWR VPWR net2151 sky130_fd_sc_hd__dlygate4sd3_1
X_06195_ net1633 _03543_ _03547_ net1207 VGND VGND VPWR VPWR _03550_ sky130_fd_sc_hd__a22o_1
Xhold511 tag_array.tag1\[3\]\[21\] VGND VGND VPWR VPWR net2162 sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 data_array.data0\[8\]\[18\] VGND VGND VPWR VPWR net2173 sky130_fd_sc_hd__dlygate4sd3_1
Xhold533 tag_array.tag1\[3\]\[24\] VGND VGND VPWR VPWR net2184 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold544 data_array.data1\[8\]\[22\] VGND VGND VPWR VPWR net2195 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold555 data_array.data1\[2\]\[9\] VGND VGND VPWR VPWR net2206 sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 tag_array.tag1\[4\]\[17\] VGND VGND VPWR VPWR net2217 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold577 data_array.data1\[14\]\[17\] VGND VGND VPWR VPWR net2228 sky130_fd_sc_hd__dlygate4sd3_1
Xhold588 data_array.data1\[8\]\[42\] VGND VGND VPWR VPWR net2239 sky130_fd_sc_hd__dlygate4sd3_1
X_09954_ net1013 net3975 net377 VGND VGND VPWR VPWR _01703_ sky130_fd_sc_hd__mux2_1
Xhold599 data_array.data0\[8\]\[46\] VGND VGND VPWR VPWR net2250 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08905_ net884 net3964 net435 VGND VGND VPWR VPWR _00662_ sky130_fd_sc_hd__mux2_1
XFILLER_103_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_46 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09885_ net929 net4252 net379 VGND VGND VPWR VPWR _01635_ sky130_fd_sc_hd__mux2_1
Xhold1200 data_array.data0\[13\]\[11\] VGND VGND VPWR VPWR net2851 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1063 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1211 tag_array.dirty1\[9\] VGND VGND VPWR VPWR net2862 sky130_fd_sc_hd__dlygate4sd3_1
X_08836_ net2018 net903 net444 VGND VGND VPWR VPWR _00594_ sky130_fd_sc_hd__mux2_1
XFILLER_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1222 lru_array.lru_mem\[2\] VGND VGND VPWR VPWR net2873 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1233 data_array.data1\[12\]\[3\] VGND VGND VPWR VPWR net2884 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1244 tag_array.tag0\[4\]\[1\] VGND VGND VPWR VPWR net2895 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1255 data_array.data0\[5\]\[22\] VGND VGND VPWR VPWR net2906 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1266 tag_array.tag1\[1\]\[12\] VGND VGND VPWR VPWR net2917 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1277 data_array.data1\[13\]\[30\] VGND VGND VPWR VPWR net2928 sky130_fd_sc_hd__dlygate4sd3_1
X_08767_ net754 net3071 net451 VGND VGND VPWR VPWR _00526_ sky130_fd_sc_hd__mux2_1
Xhold1288 tag_array.tag0\[15\]\[17\] VGND VGND VPWR VPWR net2939 sky130_fd_sc_hd__dlygate4sd3_1
X_05979_ data_array.rdata1\[49\] net832 net841 VGND VGND VPWR VPWR _03447_ sky130_fd_sc_hd__a21o_1
Xhold1299 data_array.data1\[9\]\[26\] VGND VGND VPWR VPWR net2950 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_140_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07718_ data_array.data1\[1\]\[25\] net1519 net1423 data_array.data1\[2\]\[25\] VGND
+ VGND VPWR VPWR _04934_ sky130_fd_sc_hd__a22o_1
XFILLER_25_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08698_ net2023 net730 net486 VGND VGND VPWR VPWR _00457_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07649_ _04870_ _04871_ VGND VGND VPWR VPWR _00073_ sky130_fd_sc_hd__or2_1
XFILLER_81_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10660_ net3027 net1078 net479 VGND VGND VPWR VPWR _02405_ sky130_fd_sc_hd__mux2_1
XFILLER_40_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09319_ net702 net2497 net546 VGND VGND VPWR VPWR _01073_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_114_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_114_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10591_ net2797 net1098 net471 VGND VGND VPWR VPWR _02336_ sky130_fd_sc_hd__mux2_1
X_12330_ clknet_leaf_118_clk _00003_ VGND VGND VPWR VPWR data_array.rdata0\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12261_ clknet_leaf_187_clk _01019_ VGND VGND VPWR VPWR tag_array.tag1\[14\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_14000_ clknet_leaf_123_clk _02629_ VGND VGND VPWR VPWR data_array.data1\[5\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_79_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11212_ net925 net3778 net648 VGND VGND VPWR VPWR _02955_ sky130_fd_sc_hd__mux2_1
XFILLER_181_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12192_ clknet_leaf_182_clk _01000_ VGND VGND VPWR VPWR tag_array.tag0\[14\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_122_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11143_ net947 net3233 net541 VGND VGND VPWR VPWR _02886_ sky130_fd_sc_hd__mux2_1
X_11074_ net3100 net964 net335 VGND VGND VPWR VPWR _02817_ sky130_fd_sc_hd__mux2_1
XFILLER_95_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput120 mem_rdata[29] VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_1
Xinput131 mem_rdata[39] VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10025_ net985 net2782 net561 VGND VGND VPWR VPWR _01774_ sky130_fd_sc_hd__mux2_1
Xinput142 mem_rdata[49] VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_1
Xinput153 mem_rdata[59] VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_160_3438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput164 net1694 VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__buf_2
Xhold2490 data_array.data1\[6\]\[13\] VGND VGND VPWR VPWR net4141 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11976_ clknet_leaf_25_clk _00784_ VGND VGND VPWR VPWR data_array.data0\[4\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
X_13715_ clknet_leaf_36_clk _02344_ VGND VGND VPWR VPWR data_array.data1\[1\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_10927_ net1034 net2335 net532 VGND VGND VPWR VPWR _02672_ sky130_fd_sc_hd__mux2_1
XFILLER_71_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13646_ clknet_leaf_268_clk _02275_ VGND VGND VPWR VPWR data_array.data1\[15\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10858_ net1054 net4263 net519 VGND VGND VPWR VPWR _02603_ sky130_fd_sc_hd__mux2_1
XFILLER_60_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13577_ clknet_leaf_248_clk _02206_ VGND VGND VPWR VPWR data_array.data0\[9\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_105_clk clknet_5_24__leaf_clk VGND VGND VPWR VPWR clknet_leaf_105_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_169_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10789_ net2013 net1074 net508 VGND VGND VPWR VPWR _02534_ sky130_fd_sc_hd__mux2_1
XFILLER_173_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_5_17__f_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_5_17__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_12528_ clknet_leaf_104_clk _01222_ VGND VGND VPWR VPWR tag_array.tag1\[11\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_136_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12459_ clknet_leaf_34_clk _01153_ VGND VGND VPWR VPWR data_array.data1\[9\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_10_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_184_3906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_184_3917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14129_ clknet_leaf_260_clk _02758_ VGND VGND VPWR VPWR data_array.data0\[1\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06951_ data_array.data0\[8\]\[19\] net1389 net1295 data_array.data0\[11\]\[19\]
+ _04236_ VGND VGND VPWR VPWR _04237_ sky130_fd_sc_hd__a221o_1
XFILLER_140_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05902_ net114 net1153 _03394_ _03395_ VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__a22o_1
XFILLER_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09670_ net708 net3441 net614 VGND VGND VPWR VPWR _01422_ sky130_fd_sc_hd__mux2_1
X_06882_ data_array.data0\[1\]\[13\] net1548 net1452 data_array.data0\[2\]\[13\] VGND
+ VGND VPWR VPWR _04174_ sky130_fd_sc_hd__a22o_1
X_08621_ net740 net4529 net524 VGND VGND VPWR VPWR _00380_ sky130_fd_sc_hd__mux2_1
X_05833_ net99 net1153 net1145 _03349_ VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_85_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_941 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08552_ net747 net3886 net585 VGND VGND VPWR VPWR _00320_ sky130_fd_sc_hd__mux2_1
X_05764_ _03277_ _03278_ _03279_ _03280_ VGND VGND VPWR VPWR _03281_ sky130_fd_sc_hd__or4_1
X_07503_ data_array.data1\[4\]\[5\] net1360 net1266 data_array.data1\[7\]\[5\] _04738_
+ VGND VGND VPWR VPWR _04739_ sky130_fd_sc_hd__a221o_1
X_08483_ net824 _05558_ VGND VGND VPWR VPWR _05559_ sky130_fd_sc_hd__or2_1
XFILLER_51_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05695_ _03197_ _03211_ _03206_ _03202_ VGND VGND VPWR VPWR _03212_ sky130_fd_sc_hd__or4_4
XFILLER_50_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07434_ data_array.data0\[9\]\[63\] net1548 net1452 data_array.data0\[10\]\[63\]
+ VGND VGND VPWR VPWR _04676_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_21_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07365_ data_array.data0\[12\]\[57\] net1349 net1255 data_array.data0\[15\]\[57\]
+ _04612_ VGND VGND VPWR VPWR _04613_ sky130_fd_sc_hd__a221o_1
XFILLER_148_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09104_ net869 net4216 net416 VGND VGND VPWR VPWR _00858_ sky130_fd_sc_hd__mux2_1
XFILLER_182_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06316_ net1207 _03653_ _03657_ net1633 VGND VGND VPWR VPWR _03660_ sky130_fd_sc_hd__a22o_1
XFILLER_109_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07296_ net1169 _04545_ _04549_ net1217 VGND VGND VPWR VPWR _04551_ sky130_fd_sc_hd__a22o_1
XFILLER_108_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09035_ net2003 net884 net419 VGND VGND VPWR VPWR _00790_ sky130_fd_sc_hd__mux2_1
X_06247_ tag_array.tag0\[8\]\[5\] net1410 net1316 tag_array.tag0\[11\]\[5\] _03596_
+ VGND VGND VPWR VPWR _03597_ sky130_fd_sc_hd__a221o_1
XFILLER_184_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold330 data_array.data1\[4\]\[59\] VGND VGND VPWR VPWR net1981 sky130_fd_sc_hd__dlygate4sd3_1
Xhold341 data_array.data0\[0\]\[60\] VGND VGND VPWR VPWR net1992 sky130_fd_sc_hd__dlygate4sd3_1
X_06178_ tag_array.valid1\[1\] net1557 net1461 tag_array.valid1\[2\] VGND VGND VPWR
+ VPWR _03534_ sky130_fd_sc_hd__a22o_1
XFILLER_144_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold352 data_array.data0\[4\]\[56\] VGND VGND VPWR VPWR net2003 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold363 data_array.data0\[2\]\[58\] VGND VGND VPWR VPWR net2014 sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 data_array.data1\[2\]\[27\] VGND VGND VPWR VPWR net2025 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold385 data_array.data1\[0\]\[14\] VGND VGND VPWR VPWR net2036 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 data_array.data1\[0\]\[36\] VGND VGND VPWR VPWR net2047 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout810 _05364_ VGND VGND VPWR VPWR net810 sky130_fd_sc_hd__clkbuf_2
Xfanout821 net823 VGND VGND VPWR VPWR net821 sky130_fd_sc_hd__clkbuf_2
Xfanout832 net833 VGND VGND VPWR VPWR net832 sky130_fd_sc_hd__buf_8
X_09937_ net1080 net3877 net377 VGND VGND VPWR VPWR _01686_ sky130_fd_sc_hd__mux2_1
Xfanout843 net844 VGND VGND VPWR VPWR net843 sky130_fd_sc_hd__buf_6
XFILLER_77_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout854 _05554_ VGND VGND VPWR VPWR net854 sky130_fd_sc_hd__clkbuf_2
Xfanout865 _05542_ VGND VGND VPWR VPWR net865 sky130_fd_sc_hd__buf_1
XFILLER_86_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_142_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout876 net877 VGND VGND VPWR VPWR net876 sky130_fd_sc_hd__clkbuf_2
Xfanout887 _05532_ VGND VGND VPWR VPWR net887 sky130_fd_sc_hd__buf_1
X_09868_ net998 net4619 net382 VGND VGND VPWR VPWR _01618_ sky130_fd_sc_hd__mux2_1
XFILLER_100_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1030 data_array.data0\[6\]\[16\] VGND VGND VPWR VPWR net2681 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout898 _05526_ VGND VGND VPWR VPWR net898 sky130_fd_sc_hd__clkbuf_2
XFILLER_58_565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1041 tag_array.tag0\[9\]\[10\] VGND VGND VPWR VPWR net2692 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1052 data_array.data1\[13\]\[25\] VGND VGND VPWR VPWR net2703 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08819_ net2065 net970 net443 VGND VGND VPWR VPWR _00577_ sky130_fd_sc_hd__mux2_1
Xhold1063 data_array.data0\[11\]\[42\] VGND VGND VPWR VPWR net2714 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1074 data_array.data0\[2\]\[18\] VGND VGND VPWR VPWR net2725 sky130_fd_sc_hd__dlygate4sd3_1
X_09799_ net1012 net3483 net390 VGND VGND VPWR VPWR _01550_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1085 data_array.data0\[13\]\[55\] VGND VGND VPWR VPWR net2736 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ clknet_leaf_264_clk _00638_ VGND VGND VPWR VPWR data_array.data0\[7\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1096 tag_array.tag0\[11\]\[22\] VGND VGND VPWR VPWR net2747 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_165_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11761_ clknet_leaf_229_clk _00569_ VGND VGND VPWR VPWR data_array.data0\[8\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_13500_ clknet_leaf_35_clk _02129_ VGND VGND VPWR VPWR tag_array.dirty1\[10\] sky130_fd_sc_hd__dfxtp_1
X_10712_ net2448 net870 net487 VGND VGND VPWR VPWR _02457_ sky130_fd_sc_hd__mux2_1
XFILLER_41_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14480_ clknet_leaf_172_clk _03103_ VGND VGND VPWR VPWR lru_array.lru_mem\[9\] sky130_fd_sc_hd__dfxtp_1
X_11692_ clknet_leaf_136_clk _00500_ VGND VGND VPWR VPWR tag_array.tag1\[15\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_41_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13431_ clknet_leaf_5_clk _02061_ VGND VGND VPWR VPWR data_array.data1\[8\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10643_ net2476 net890 net467 VGND VGND VPWR VPWR _02388_ sky130_fd_sc_hd__mux2_1
XFILLER_158_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13362_ clknet_leaf_142_clk _01992_ VGND VGND VPWR VPWR tag_array.tag0\[2\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_158_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10574_ net911 net4253 net453 VGND VGND VPWR VPWR _02319_ sky130_fd_sc_hd__mux2_1
XFILLER_155_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_153_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12313_ clknet_leaf_232_clk _01071_ VGND VGND VPWR VPWR tag_array.tag1\[12\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_127_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13293_ clknet_leaf_248_clk _01923_ VGND VGND VPWR VPWR data_array.data0\[10\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_114_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12244_ clknet_leaf_167_clk _01002_ VGND VGND VPWR VPWR tag_array.tag1\[14\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_108_773 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12175_ clknet_leaf_158_clk _00983_ VGND VGND VPWR VPWR tag_array.tag0\[14\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_131_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11126_ net1015 net3568 net550 VGND VGND VPWR VPWR _02869_ sky130_fd_sc_hd__mux2_1
XFILLER_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11057_ net2230 net1032 net333 VGND VGND VPWR VPWR _02800_ sky130_fd_sc_hd__mux2_1
XFILLER_114_1042 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10008_ net1054 net3239 net561 VGND VGND VPWR VPWR _01757_ sky130_fd_sc_hd__mux2_1
XFILLER_37_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_177_3754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11959_ clknet_leaf_91_clk _00767_ VGND VGND VPWR VPWR data_array.data0\[4\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_178_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_177_3765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13629_ clknet_leaf_219_clk _02258_ VGND VGND VPWR VPWR data_array.data0\[9\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_15_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07150_ data_array.data0\[5\]\[37\] net1546 net1450 data_array.data0\[6\]\[37\] VGND
+ VGND VPWR VPWR _04418_ sky130_fd_sc_hd__a22o_1
X_06101_ data_array.rdata0\[16\] net1136 net1117 data_array.rdata1\[16\] VGND VGND
+ VPWR VPWR net270 sky130_fd_sc_hd__a22o_1
X_07081_ data_array.data0\[4\]\[31\] net1384 net1290 data_array.data0\[7\]\[31\] _04354_
+ VGND VGND VPWR VPWR _04355_ sky130_fd_sc_hd__a221o_1
XFILLER_172_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06032_ net1160 net1137 net1118 net27 VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__o31a_1
XFILLER_160_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07983_ data_array.data1\[0\]\[49\] net1381 net1287 data_array.data1\[3\]\[49\] _05174_
+ VGND VGND VPWR VPWR _05175_ sky130_fd_sc_hd__a221o_1
XFILLER_87_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09722_ net698 net3515 net610 VGND VGND VPWR VPWR _01474_ sky130_fd_sc_hd__mux2_1
X_06934_ _04220_ _04221_ VGND VGND VPWR VPWR _00008_ sky130_fd_sc_hd__or2_1
XFILLER_80_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_52_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_52_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09653_ net777 net4111 net612 VGND VGND VPWR VPWR _01405_ sky130_fd_sc_hd__mux2_1
X_06865_ data_array.data0\[4\]\[11\] net1383 net1289 data_array.data0\[7\]\[11\] _04158_
+ VGND VGND VPWR VPWR _04159_ sky130_fd_sc_hd__a221o_1
XFILLER_110_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08604_ net706 net3771 net537 VGND VGND VPWR VPWR _00363_ sky130_fd_sc_hd__mux2_1
X_05816_ _03320_ _03326_ _03327_ _03332_ VGND VGND VPWR VPWR _03333_ sky130_fd_sc_hd__nor4_4
X_09584_ net1012 net3234 net398 VGND VGND VPWR VPWR _01336_ sky130_fd_sc_hd__mux2_1
X_06796_ data_array.data0\[13\]\[5\] net1550 net1454 data_array.data0\[14\]\[5\] VGND
+ VGND VPWR VPWR _04096_ sky130_fd_sc_hd__a22o_1
XFILLER_63_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_118_Right_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08535_ net813 _05561_ VGND VGND VPWR VPWR _05594_ sky130_fd_sc_hd__nand2_2
X_05747_ fsm.tag_out1\[7\] net6 VGND VGND VPWR VPWR _03264_ sky130_fd_sc_hd__and2b_1
XFILLER_35_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08466_ _03507_ _03511_ VGND VGND VPWR VPWR _05547_ sky130_fd_sc_hd__nor2_1
X_05678_ net5 fsm.tag_out0\[6\] VGND VGND VPWR VPWR _03195_ sky130_fd_sc_hd__and2b_1
XFILLER_23_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07417_ net1219 _04655_ _04659_ net1171 VGND VGND VPWR VPWR _04661_ sky130_fd_sc_hd__a22o_1
X_08397_ net134 net69 net1642 VGND VGND VPWR VPWR _05501_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_98_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07348_ data_array.data0\[5\]\[55\] net1534 net1438 data_array.data0\[6\]\[55\] VGND
+ VGND VPWR VPWR _04598_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_98_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_857 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07279_ data_array.data0\[0\]\[49\] net1380 net1286 data_array.data0\[3\]\[49\] _04534_
+ VGND VGND VPWR VPWR _04535_ sky130_fd_sc_hd__a221o_1
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09018_ net3270 net954 net421 VGND VGND VPWR VPWR _00773_ sky130_fd_sc_hd__mux2_1
XFILLER_164_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10290_ net2109 net1000 net634 VGND VGND VPWR VPWR _02037_ sky130_fd_sc_hd__mux2_1
XFILLER_145_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold160 data_array.data1\[2\]\[11\] VGND VGND VPWR VPWR net1811 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold171 tag_array.tag1\[8\]\[2\] VGND VGND VPWR VPWR net1822 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_176_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold182 data_array.data1\[1\]\[17\] VGND VGND VPWR VPWR net1833 sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 tag_array.tag1\[0\]\[1\] VGND VGND VPWR VPWR net1844 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout1605 net1606 VGND VGND VPWR VPWR net1605 sky130_fd_sc_hd__clkbuf_4
Xfanout1616 net1617 VGND VGND VPWR VPWR net1616 sky130_fd_sc_hd__buf_4
XFILLER_78_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1627 _03506_ VGND VGND VPWR VPWR net1627 sky130_fd_sc_hd__clkbuf_4
XFILLER_132_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout640 net644 VGND VGND VPWR VPWR net640 sky130_fd_sc_hd__buf_4
Xfanout1638 net1639 VGND VGND VPWR VPWR net1638 sky130_fd_sc_hd__buf_4
Xfanout1649 net163 VGND VGND VPWR VPWR net1649 sky130_fd_sc_hd__buf_2
Xfanout651 _05551_ VGND VGND VPWR VPWR net651 sky130_fd_sc_hd__clkbuf_4
Xfanout662 net666 VGND VGND VPWR VPWR net662 sky130_fd_sc_hd__buf_2
XFILLER_144_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13980_ clknet_leaf_123_clk _02609_ VGND VGND VPWR VPWR data_array.data1\[5\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout673 net676 VGND VGND VPWR VPWR net673 sky130_fd_sc_hd__buf_4
Xfanout684 net685 VGND VGND VPWR VPWR net684 sky130_fd_sc_hd__buf_4
Xfanout695 net697 VGND VGND VPWR VPWR net695 sky130_fd_sc_hd__clkbuf_2
XFILLER_46_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12931_ clknet_leaf_242_clk _01625_ VGND VGND VPWR VPWR data_array.data0\[13\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_86_682 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12862_ clknet_leaf_71_clk _01556_ VGND VGND VPWR VPWR data_array.data0\[12\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_73_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11813_ clknet_leaf_63_clk _00621_ VGND VGND VPWR VPWR data_array.data0\[7\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12793_ clknet_leaf_33_clk _01487_ VGND VGND VPWR VPWR tag_array.tag1\[10\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11744_ clknet_leaf_111_clk _00552_ VGND VGND VPWR VPWR data_array.data0\[8\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_3337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_155_3348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14463_ clknet_leaf_78_clk _03086_ VGND VGND VPWR VPWR data_array.data1\[7\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
X_11675_ clknet_leaf_139_clk _00483_ VGND VGND VPWR VPWR tag_array.tag1\[1\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_12_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_172_3662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13414_ clknet_leaf_6_clk _02044_ VGND VGND VPWR VPWR data_array.data1\[8\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_172_3673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10626_ net2095 net957 net473 VGND VGND VPWR VPWR _02371_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_116_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14394_ clknet_leaf_79_clk _03017_ VGND VGND VPWR VPWR data_array.data1\[10\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13345_ clknet_leaf_219_clk _01975_ VGND VGND VPWR VPWR data_array.data0\[10\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_133_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10557_ net978 net3869 net461 VGND VGND VPWR VPWR _02302_ sky130_fd_sc_hd__mux2_1
XFILLER_6_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13276_ clknet_leaf_61_clk _01906_ VGND VGND VPWR VPWR data_array.data0\[11\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
X_10488_ net992 net3217 net349 VGND VGND VPWR VPWR _02233_ sky130_fd_sc_hd__mux2_1
XFILLER_154_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12227_ clknet_leaf_148_clk _00180_ VGND VGND VPWR VPWR fsm.tag_out1\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_142_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12158_ clknet_leaf_163_clk _00966_ VGND VGND VPWR VPWR tag_array.tag0\[13\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_69_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11109_ net1083 net2618 net550 VGND VGND VPWR VPWR _02852_ sky130_fd_sc_hd__mux2_1
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12089_ clknet_leaf_259_clk _00897_ VGND VGND VPWR VPWR data_array.data1\[14\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_179_3805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06650_ tag_array.tag1\[12\]\[17\] net1421 net1327 tag_array.tag1\[15\]\[17\] _03962_
+ VGND VGND VPWR VPWR _03963_ sky130_fd_sc_hd__a221o_1
XFILLER_40_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06581_ net1229 _03895_ _03899_ net1181 VGND VGND VPWR VPWR _03901_ sky130_fd_sc_hd__a22o_1
X_08320_ net1127 _05449_ VGND VGND VPWR VPWR _05450_ sky130_fd_sc_hd__and2_1
XFILLER_177_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08251_ net1650 net1161 net19 VGND VGND VPWR VPWR _05402_ sky130_fd_sc_hd__and3_1
X_07202_ data_array.data0\[4\]\[42\] net1388 net1294 data_array.data0\[7\]\[42\] _04464_
+ VGND VGND VPWR VPWR _04465_ sky130_fd_sc_hd__a221o_1
X_08182_ _03146_ net827 net826 net229 VGND VGND VPWR VPWR _05353_ sky130_fd_sc_hd__o31ai_2
XFILLER_119_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07133_ data_array.data0\[9\]\[36\] net1604 net1508 data_array.data0\[10\]\[36\]
+ VGND VGND VPWR VPWR _04402_ sky130_fd_sc_hd__a22o_1
XFILLER_146_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07064_ net1202 _04333_ _04337_ net1628 VGND VGND VPWR VPWR _04340_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput210 net210 VGND VGND VPWR VPWR cpu_rdata[50] sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_93_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput221 net221 VGND VGND VPWR VPWR cpu_rdata[60] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_93_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06015_ data_array.rdata1\[61\] net831 net839 VGND VGND VPWR VPWR _03471_ sky130_fd_sc_hd__a21o_1
Xoutput232 net232 VGND VGND VPWR VPWR mem_addr[11] sky130_fd_sc_hd__buf_2
Xoutput243 net243 VGND VGND VPWR VPWR mem_addr[21] sky130_fd_sc_hd__buf_2
Xoutput254 net254 VGND VGND VPWR VPWR mem_addr[31] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput265 net265 VGND VGND VPWR VPWR mem_wdata[11] sky130_fd_sc_hd__buf_2
XFILLER_99_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput276 net276 VGND VGND VPWR VPWR mem_wdata[21] sky130_fd_sc_hd__buf_2
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput287 net287 VGND VGND VPWR VPWR mem_wdata[31] sky130_fd_sc_hd__buf_2
Xoutput298 net298 VGND VGND VPWR VPWR mem_wdata[41] sky130_fd_sc_hd__buf_2
XFILLER_102_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07966_ net1632 _05153_ _05157_ net1206 VGND VGND VPWR VPWR _05160_ sky130_fd_sc_hd__a22o_1
X_09705_ net768 net2688 net609 VGND VGND VPWR VPWR _01457_ sky130_fd_sc_hd__mux2_1
X_06917_ data_array.data0\[13\]\[16\] net1549 net1453 data_array.data0\[14\]\[16\]
+ VGND VGND VPWR VPWR _04206_ sky130_fd_sc_hd__a22o_1
X_07897_ data_array.data1\[12\]\[41\] net1336 net1242 data_array.data1\[15\]\[41\]
+ _05096_ VGND VGND VPWR VPWR _05097_ sky130_fd_sc_hd__a221o_1
XFILLER_74_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_94_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_94_clk sky130_fd_sc_hd__clkbuf_8
X_09636_ net744 net3141 net615 VGND VGND VPWR VPWR _01388_ sky130_fd_sc_hd__mux2_1
X_06848_ data_array.data0\[8\]\[10\] net1411 net1317 data_array.data0\[11\]\[10\]
+ _04142_ VGND VGND VPWR VPWR _04143_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09567_ net1080 net3205 net400 VGND VGND VPWR VPWR _01319_ sky130_fd_sc_hd__mux2_1
X_06779_ net1176 _04075_ _04079_ net1224 VGND VGND VPWR VPWR _04081_ sky130_fd_sc_hd__a22o_1
XFILLER_82_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08518_ _03516_ _03519_ VGND VGND VPWR VPWR _05583_ sky130_fd_sc_hd__nor2_2
XFILLER_130_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09498_ net736 net2289 net624 VGND VGND VPWR VPWR _01251_ sky130_fd_sc_hd__mux2_1
X_08449_ net1126 _05535_ VGND VGND VPWR VPWR _05536_ sky130_fd_sc_hd__and2_1
XFILLER_12_958 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11460_ clknet_leaf_53_clk _00270_ VGND VGND VPWR VPWR data_array.data0\[0\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_109_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10411_ net2716 net1008 net661 VGND VGND VPWR VPWR _02157_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_150_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11391_ clknet_leaf_133_clk _00201_ VGND VGND VPWR VPWR tag_array.tag1\[7\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_150_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_1025 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13130_ clknet_leaf_108_clk _01824_ VGND VGND VPWR VPWR tag_array.tag0\[3\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_10342_ net732 net3573 net591 VGND VGND VPWR VPWR _02089_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13061_ clknet_leaf_85_clk _01755_ VGND VGND VPWR VPWR data_array.data1\[13\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_10273_ net1982 net1070 net640 VGND VGND VPWR VPWR _02020_ sky130_fd_sc_hd__mux2_1
XFILLER_3_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12012_ clknet_leaf_9_clk _00820_ VGND VGND VPWR VPWR data_array.data0\[6\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1402 net1403 VGND VGND VPWR VPWR net1402 sky130_fd_sc_hd__clkbuf_4
XFILLER_120_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1413 net1422 VGND VGND VPWR VPWR net1413 sky130_fd_sc_hd__clkbuf_4
Xfanout1424 net1425 VGND VGND VPWR VPWR net1424 sky130_fd_sc_hd__clkbuf_4
Xfanout1435 net1437 VGND VGND VPWR VPWR net1435 sky130_fd_sc_hd__clkbuf_4
Xfanout1446 net1447 VGND VGND VPWR VPWR net1446 sky130_fd_sc_hd__buf_2
Xfanout1457 net1458 VGND VGND VPWR VPWR net1457 sky130_fd_sc_hd__clkbuf_4
Xfanout470 net477 VGND VGND VPWR VPWR net470 sky130_fd_sc_hd__clkbuf_8
Xfanout1468 net1470 VGND VGND VPWR VPWR net1468 sky130_fd_sc_hd__clkbuf_4
Xfanout481 net482 VGND VGND VPWR VPWR net481 sky130_fd_sc_hd__buf_4
XFILLER_48_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1479 net1480 VGND VGND VPWR VPWR net1479 sky130_fd_sc_hd__clkbuf_4
Xfanout492 net495 VGND VGND VPWR VPWR net492 sky130_fd_sc_hd__clkbuf_8
X_13963_ clknet_leaf_28_clk _02592_ VGND VGND VPWR VPWR data_array.data1\[5\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_109_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_85_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_85_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_58_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12914_ clknet_leaf_15_clk _01608_ VGND VGND VPWR VPWR data_array.data0\[13\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_13894_ clknet_leaf_120_clk _02523_ VGND VGND VPWR VPWR data_array.data1\[3\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12845_ clknet_leaf_192_clk _01539_ VGND VGND VPWR VPWR data_array.data0\[12\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_174_3702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12776_ clknet_leaf_106_clk _01470_ VGND VGND VPWR VPWR tag_array.tag0\[6\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_159_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11727_ clknet_leaf_185_clk _00535_ VGND VGND VPWR VPWR tag_array.tag0\[9\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_148_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14446_ clknet_leaf_69_clk _03069_ VGND VGND VPWR VPWR data_array.data1\[7\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_11658_ clknet_leaf_189_clk _00466_ VGND VGND VPWR VPWR tag_array.tag1\[2\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_80_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_980 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10609_ net2325 net1025 net470 VGND VGND VPWR VPWR _02354_ sky130_fd_sc_hd__mux2_1
XFILLER_128_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14377_ clknet_leaf_248_clk _03000_ VGND VGND VPWR VPWR data_array.data1\[10\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_11589_ clknet_leaf_135_clk _00397_ VGND VGND VPWR VPWR tag_array.tag1\[4\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_127_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold907 data_array.data1\[6\]\[16\] VGND VGND VPWR VPWR net2558 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13328_ clknet_leaf_218_clk _01958_ VGND VGND VPWR VPWR data_array.data0\[10\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold918 data_array.data1\[13\]\[54\] VGND VGND VPWR VPWR net2569 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_170_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold929 data_array.data0\[4\]\[21\] VGND VGND VPWR VPWR net2580 sky130_fd_sc_hd__dlygate4sd3_1
X_13259_ clknet_leaf_260_clk _01889_ VGND VGND VPWR VPWR data_array.data0\[11\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_143_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2308 data_array.data0\[3\]\[22\] VGND VGND VPWR VPWR net3959 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2319 data_array.data1\[15\]\[25\] VGND VGND VPWR VPWR net3970 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07820_ data_array.data1\[8\]\[34\] net1341 net1247 data_array.data1\[11\]\[34\]
+ _05026_ VGND VGND VPWR VPWR _05027_ sky130_fd_sc_hd__a221o_1
Xhold1607 data_array.data1\[6\]\[27\] VGND VGND VPWR VPWR net3258 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1618 tag_array.tag0\[10\]\[16\] VGND VGND VPWR VPWR net3269 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1629 data_array.data1\[11\]\[13\] VGND VGND VPWR VPWR net3280 sky130_fd_sc_hd__dlygate4sd3_1
X_07751_ data_array.data1\[5\]\[28\] net1540 net1444 data_array.data1\[6\]\[28\] VGND
+ VGND VPWR VPWR _04964_ sky130_fd_sc_hd__a22o_1
XFILLER_37_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_76_clk clknet_5_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_76_clk sky130_fd_sc_hd__clkbuf_8
X_06702_ net1182 _04005_ _04009_ net1230 VGND VGND VPWR VPWR _04011_ sky130_fd_sc_hd__a22o_1
X_07682_ _04900_ _04901_ VGND VGND VPWR VPWR _00077_ sky130_fd_sc_hd__or2_1
XFILLER_25_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09421_ net980 net3306 net578 VGND VGND VPWR VPWR _01174_ sky130_fd_sc_hd__mux2_1
XFILLER_92_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_622 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06633_ tag_array.tag1\[5\]\[15\] net1575 net1479 tag_array.tag1\[6\]\[15\] VGND
+ VGND VPWR VPWR _03948_ sky130_fd_sc_hd__a22o_1
XFILLER_53_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09352_ net993 net3391 net407 VGND VGND VPWR VPWR _01105_ sky130_fd_sc_hd__mux2_1
X_06564_ tag_array.tag1\[4\]\[9\] net1418 net1324 tag_array.tag1\[7\]\[9\] _03884_
+ VGND VGND VPWR VPWR _03885_ sky130_fd_sc_hd__a221o_1
XFILLER_166_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08303_ net1782 net1072 net691 VGND VGND VPWR VPWR _00230_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09283_ net746 net3350 net563 VGND VGND VPWR VPWR _01037_ sky130_fd_sc_hd__mux2_1
XFILLER_127_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06495_ tag_array.tag1\[9\]\[3\] net1561 net1465 tag_array.tag1\[10\]\[3\] VGND VGND
+ VPWR VPWR _03822_ sky130_fd_sc_hd__a22o_1
X_08234_ fsm.tag_out1\[13\] net818 net810 fsm.tag_out0\[13\] _05390_ VGND VGND VPWR
+ VPWR _05391_ sky130_fd_sc_hd__a221o_2
XFILLER_138_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08165_ net1230 _05335_ _05339_ net1182 VGND VGND VPWR VPWR _05341_ sky130_fd_sc_hd__a22o_1
X_07116_ data_array.data0\[8\]\[34\] net1340 net1246 data_array.data0\[11\]\[34\]
+ _04386_ VGND VGND VPWR VPWR _04387_ sky130_fd_sc_hd__a221o_1
XFILLER_180_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08096_ data_array.data1\[5\]\[59\] net1570 net1474 data_array.data1\[6\]\[59\] VGND
+ VGND VPWR VPWR _05278_ sky130_fd_sc_hd__a22o_1
XFILLER_118_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload80 clknet_leaf_54_clk VGND VGND VPWR VPWR clkload80/Y sky130_fd_sc_hd__bufinv_16
Xclkload91 clknet_leaf_64_clk VGND VGND VPWR VPWR clkload91/Y sky130_fd_sc_hd__clkinvlp_4
X_07047_ data_array.data0\[5\]\[28\] net1540 net1444 data_array.data0\[6\]\[28\] VGND
+ VGND VPWR VPWR _04324_ sky130_fd_sc_hd__a22o_1
XFILLER_0_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_12 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2820 data_array.data1\[3\]\[42\] VGND VGND VPWR VPWR net4471 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2831 data_array.data1\[11\]\[6\] VGND VGND VPWR VPWR net4482 sky130_fd_sc_hd__dlygate4sd3_1
X_08998_ net1803 net1032 net422 VGND VGND VPWR VPWR _00753_ sky130_fd_sc_hd__mux2_1
Xhold2842 data_array.data1\[15\]\[53\] VGND VGND VPWR VPWR net4493 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2853 data_array.data1\[5\]\[59\] VGND VGND VPWR VPWR net4504 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2864 data_array.data0\[11\]\[55\] VGND VGND VPWR VPWR net4515 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2875 data_array.data0\[11\]\[56\] VGND VGND VPWR VPWR net4526 sky130_fd_sc_hd__dlygate4sd3_1
X_07949_ data_array.data1\[5\]\[46\] net1524 net1428 data_array.data1\[6\]\[46\] VGND
+ VGND VPWR VPWR _05144_ sky130_fd_sc_hd__a22o_1
Xhold2886 tag_array.tag0\[5\]\[9\] VGND VGND VPWR VPWR net4537 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_67_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_67_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_28_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2897 data_array.data1\[7\]\[11\] VGND VGND VPWR VPWR net4548 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_170_Right_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10960_ net900 net3833 net528 VGND VGND VPWR VPWR _02705_ sky130_fd_sc_hd__mux2_1
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09619_ net873 net3981 net398 VGND VGND VPWR VPWR _01371_ sky130_fd_sc_hd__mux2_1
X_10891_ _05514_ net2523 net521 VGND VGND VPWR VPWR _02636_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12630_ clknet_leaf_104_clk _01324_ VGND VGND VPWR VPWR data_array.data0\[15\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_43_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_84_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12561_ clknet_leaf_182_clk _01255_ VGND VGND VPWR VPWR tag_array.tag0\[11\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_14300_ clknet_leaf_131_clk _02929_ VGND VGND VPWR VPWR data_array.data1\[11\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_11512_ clknet_leaf_33_clk _00320_ VGND VGND VPWR VPWR tag_array.tag1\[9\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_141_1027 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12492_ clknet_leaf_80_clk _01186_ VGND VGND VPWR VPWR data_array.data1\[9\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_156_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14231_ clknet_leaf_70_clk _02860_ VGND VGND VPWR VPWR data_array.data1\[12\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_11443_ clknet_leaf_260_clk _00253_ VGND VGND VPWR VPWR data_array.data0\[0\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14162_ clknet_leaf_112_clk _02791_ VGND VGND VPWR VPWR data_array.data0\[2\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_11374_ net1647 net2420 net631 VGND VGND VPWR VPWR _03117_ sky130_fd_sc_hd__mux2_1
XFILLER_152_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13113_ clknet_leaf_106_clk _01807_ VGND VGND VPWR VPWR tag_array.tag0\[3\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_124_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10325_ net1869 net862 net642 VGND VGND VPWR VPWR _02072_ sky130_fd_sc_hd__mux2_1
X_14093_ clknet_leaf_209_clk _02722_ VGND VGND VPWR VPWR data_array.data0\[1\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_180_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13044_ clknet_leaf_51_clk _01738_ VGND VGND VPWR VPWR data_array.data0\[3\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
X_10256_ net721 net2774 net598 VGND VGND VPWR VPWR _02003_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_167_3572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1210 net1211 VGND VGND VPWR VPWR net1210 sky130_fd_sc_hd__buf_4
XFILLER_79_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1221 net1222 VGND VGND VPWR VPWR net1221 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_128_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1232 net1233 VGND VGND VPWR VPWR net1232 sky130_fd_sc_hd__clkbuf_4
X_10187_ net1059 net3263 net356 VGND VGND VPWR VPWR _01934_ sky130_fd_sc_hd__mux2_1
Xfanout1243 net1244 VGND VGND VPWR VPWR net1243 sky130_fd_sc_hd__clkbuf_4
XFILLER_78_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_128_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1254 net1258 VGND VGND VPWR VPWR net1254 sky130_fd_sc_hd__buf_2
Xfanout1265 net1266 VGND VGND VPWR VPWR net1265 sky130_fd_sc_hd__clkbuf_4
XFILLER_93_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1276 net1282 VGND VGND VPWR VPWR net1276 sky130_fd_sc_hd__buf_2
Xfanout1287 net1288 VGND VGND VPWR VPWR net1287 sky130_fd_sc_hd__clkbuf_4
XFILLER_8_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_58_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_58_clk sky130_fd_sc_hd__clkbuf_8
Xfanout1298 net1306 VGND VGND VPWR VPWR net1298 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_4_11_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_11_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_93_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13946_ clknet_leaf_246_clk _02575_ VGND VGND VPWR VPWR data_array.data1\[4\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_335 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13877_ clknet_leaf_26_clk _02506_ VGND VGND VPWR VPWR data_array.data1\[3\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_179_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12828_ clknet_leaf_101_clk _01522_ VGND VGND VPWR VPWR tag_array.tag1\[0\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_12759_ clknet_leaf_168_clk _01453_ VGND VGND VPWR VPWR tag_array.tag0\[6\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_06280_ tag_array.tag0\[12\]\[8\] net1410 net1316 tag_array.tag0\[15\]\[8\] _03626_
+ VGND VGND VPWR VPWR _03627_ sky130_fd_sc_hd__a221o_1
X_14429_ clknet_leaf_200_clk _03052_ VGND VGND VPWR VPWR data_array.data1\[7\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_42_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold704 tag_array.tag0\[13\]\[2\] VGND VGND VPWR VPWR net2355 sky130_fd_sc_hd__dlygate4sd3_1
Xhold715 data_array.data0\[14\]\[56\] VGND VGND VPWR VPWR net2366 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_944 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold726 tag_array.tag1\[4\]\[6\] VGND VGND VPWR VPWR net2377 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold737 data_array.data0\[1\]\[12\] VGND VGND VPWR VPWR net2388 sky130_fd_sc_hd__dlygate4sd3_1
X_09970_ net948 net2970 net377 VGND VGND VPWR VPWR _01719_ sky130_fd_sc_hd__mux2_1
Xhold748 data_array.data0\[1\]\[28\] VGND VGND VPWR VPWR net2399 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold759 data_array.data0\[0\]\[58\] VGND VGND VPWR VPWR net2410 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08921_ net1080 net2821 net432 VGND VGND VPWR VPWR _00677_ sky130_fd_sc_hd__mux2_1
XFILLER_131_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2105 data_array.data0\[7\]\[44\] VGND VGND VPWR VPWR net3756 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2116 data_array.data1\[6\]\[41\] VGND VGND VPWR VPWR net3767 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2127 data_array.data1\[11\]\[46\] VGND VGND VPWR VPWR net3778 sky130_fd_sc_hd__dlygate4sd3_1
X_08852_ net1096 net3977 net439 VGND VGND VPWR VPWR _00609_ sky130_fd_sc_hd__mux2_1
Xhold2138 data_array.data0\[15\]\[37\] VGND VGND VPWR VPWR net3789 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2149 data_array.data0\[11\]\[38\] VGND VGND VPWR VPWR net3800 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1404 tag_array.tag0\[1\]\[12\] VGND VGND VPWR VPWR net3055 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1415 data_array.data0\[11\]\[13\] VGND VGND VPWR VPWR net3066 sky130_fd_sc_hd__dlygate4sd3_1
X_07803_ _05010_ _05011_ VGND VGND VPWR VPWR _00089_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_179_Left_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1426 data_array.data1\[5\]\[23\] VGND VGND VPWR VPWR net3077 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1437 data_array.data1\[12\]\[27\] VGND VGND VPWR VPWR net3088 sky130_fd_sc_hd__dlygate4sd3_1
X_08783_ net807 _05556_ VGND VGND VPWR VPWR _05607_ sky130_fd_sc_hd__and2_1
X_05995_ net148 net1152 _03456_ _03457_ VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__a22o_1
Xhold1448 tag_array.tag0\[3\]\[13\] VGND VGND VPWR VPWR net3099 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_88_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_49_clk clknet_5_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_49_clk sky130_fd_sc_hd__clkbuf_8
Xhold1459 data_array.data1\[11\]\[14\] VGND VGND VPWR VPWR net3110 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_88_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07734_ data_array.data1\[0\]\[26\] net1335 net1241 data_array.data1\[3\]\[26\] _04948_
+ VGND VGND VPWR VPWR _04949_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_0_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07665_ data_array.data1\[9\]\[20\] net1610 net1514 data_array.data1\[10\]\[20\]
+ VGND VGND VPWR VPWR _04886_ sky130_fd_sc_hd__a22o_1
XFILLER_26_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09404_ net1050 net3760 net586 VGND VGND VPWR VPWR _01157_ sky130_fd_sc_hd__mux2_1
X_06616_ tag_array.tag1\[9\]\[14\] net1558 net1462 tag_array.tag1\[10\]\[14\] VGND
+ VGND VPWR VPWR _03932_ sky130_fd_sc_hd__a22o_1
XFILLER_80_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07596_ data_array.data1\[8\]\[14\] net1378 net1284 data_array.data1\[11\]\[14\]
+ _04822_ VGND VGND VPWR VPWR _04823_ sky130_fd_sc_hd__a221o_1
XFILLER_164_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09335_ net1061 net3952 net408 VGND VGND VPWR VPWR _01088_ sky130_fd_sc_hd__mux2_1
X_06547_ net1636 _03863_ _03867_ net1210 VGND VGND VPWR VPWR _03870_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_62_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09266_ net714 net3947 net573 VGND VGND VPWR VPWR _01020_ sky130_fd_sc_hd__mux2_1
X_06478_ tag_array.tag1\[8\]\[1\] net1368 net1274 tag_array.tag1\[11\]\[1\] _03806_
+ VGND VGND VPWR VPWR _03807_ sky130_fd_sc_hd__a221o_1
X_08217_ net764 net3980 net804 VGND VGND VPWR VPWR _00203_ sky130_fd_sc_hd__mux2_1
XFILLER_166_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09197_ net794 net2451 net631 VGND VGND VPWR VPWR _00951_ sky130_fd_sc_hd__mux2_1
XFILLER_101_1022 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08148_ tag_array.dirty1\[0\] net1350 net1256 tag_array.dirty1\[3\] _05324_ VGND
+ VGND VPWR VPWR _05325_ sky130_fd_sc_hd__a221o_1
XFILLER_136_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08079_ data_array.data1\[9\]\[58\] net1551 net1455 data_array.data1\[10\]\[58\]
+ VGND VGND VPWR VPWR _05262_ sky130_fd_sc_hd__a22o_1
Xclkload180 clknet_leaf_180_clk VGND VGND VPWR VPWR clkload180/Y sky130_fd_sc_hd__inv_8
Xclkload191 clknet_leaf_100_clk VGND VGND VPWR VPWR clkload191/Y sky130_fd_sc_hd__clkinv_2
XFILLER_162_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10110_ net1105 net4384 net362 VGND VGND VPWR VPWR _01858_ sky130_fd_sc_hd__mux2_1
X_11090_ net2860 net903 net330 VGND VGND VPWR VPWR _02833_ sky130_fd_sc_hd__mux2_1
XFILLER_0_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10041_ net923 net3989 net563 VGND VGND VPWR VPWR _01790_ sky130_fd_sc_hd__mux2_1
XFILLER_0_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_145_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_145_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2650 data_array.data0\[15\]\[4\] VGND VGND VPWR VPWR net4301 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 tag_array.valid0\[14\] VGND VGND VPWR VPWR net1704 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2661 tag_array.dirty0\[6\] VGND VGND VPWR VPWR net4312 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2672 data_array.data1\[7\]\[7\] VGND VGND VPWR VPWR net4323 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 tag_array.valid0\[15\] VGND VGND VPWR VPWR net1715 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2683 data_array.data1\[15\]\[57\] VGND VGND VPWR VPWR net4334 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2694 data_array.data1\[13\]\[38\] VGND VGND VPWR VPWR net4345 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_162_3480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold75 tag_array.tag1\[2\]\[18\] VGND VGND VPWR VPWR net1726 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold86 data_array.data0\[4\]\[15\] VGND VGND VPWR VPWR net1737 sky130_fd_sc_hd__dlygate4sd3_1
X_13800_ clknet_leaf_257_clk _02429_ VGND VGND VPWR VPWR data_array.data1\[2\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1960 tag_array.tag1\[12\]\[24\] VGND VGND VPWR VPWR net3611 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 data_array.data1\[1\]\[44\] VGND VGND VPWR VPWR net1748 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1971 data_array.data0\[3\]\[20\] VGND VGND VPWR VPWR net3622 sky130_fd_sc_hd__dlygate4sd3_1
X_11992_ clknet_leaf_247_clk _00800_ VGND VGND VPWR VPWR data_array.data0\[6\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_57_983 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1982 tag_array.tag1\[13\]\[2\] VGND VGND VPWR VPWR net3633 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1993 data_array.data0\[9\]\[59\] VGND VGND VPWR VPWR net3644 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_123_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13731_ clknet_leaf_248_clk _02360_ VGND VGND VPWR VPWR data_array.data1\[1\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_10943_ net968 net3873 net527 VGND VGND VPWR VPWR _02688_ sky130_fd_sc_hd__mux2_1
XFILLER_21_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10874_ net990 net2902 net520 VGND VGND VPWR VPWR _02619_ sky130_fd_sc_hd__mux2_1
X_13662_ clknet_leaf_24_clk _02291_ VGND VGND VPWR VPWR data_array.data1\[15\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_43_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12613_ clknet_leaf_168_clk _01307_ VGND VGND VPWR VPWR tag_array.tag0\[0\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_13593_ clknet_leaf_48_clk _02222_ VGND VGND VPWR VPWR data_array.data0\[9\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_169_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12544_ clknet_leaf_164_clk _01238_ VGND VGND VPWR VPWR tag_array.tag0\[11\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12475_ clknet_leaf_248_clk _01169_ VGND VGND VPWR VPWR data_array.data1\[9\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_169_3601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11426_ clknet_leaf_63_clk _00236_ VGND VGND VPWR VPWR data_array.data0\[0\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_14214_ clknet_leaf_111_clk _02843_ VGND VGND VPWR VPWR data_array.data0\[2\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_169_3612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_6 _00119_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14145_ clknet_leaf_234_clk _02774_ VGND VGND VPWR VPWR data_array.data0\[1\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
X_11357_ net864 net3168 net799 VGND VGND VPWR VPWR _03100_ sky130_fd_sc_hd__mux2_1
XFILLER_152_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10308_ net1800 net931 net635 VGND VGND VPWR VPWR _02055_ sky130_fd_sc_hd__mux2_1
XFILLER_152_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14076_ clknet_leaf_212_clk _02705_ VGND VGND VPWR VPWR data_array.data1\[6\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
X_11288_ net879 net3512 net677 VGND VGND VPWR VPWR _03031_ sky130_fd_sc_hd__mux2_1
XFILLER_79_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13027_ clknet_leaf_93_clk _01721_ VGND VGND VPWR VPWR data_array.data0\[3\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
X_10239_ net788 net2856 net595 VGND VGND VPWR VPWR _01986_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_182_3856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1051 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1040 _05454_ VGND VGND VPWR VPWR net1040 sky130_fd_sc_hd__clkbuf_2
Xfanout1051 _05450_ VGND VGND VPWR VPWR net1051 sky130_fd_sc_hd__clkbuf_2
Xfanout1062 _05444_ VGND VGND VPWR VPWR net1062 sky130_fd_sc_hd__clkbuf_2
XFILLER_66_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1073 _05438_ VGND VGND VPWR VPWR net1073 sky130_fd_sc_hd__buf_1
Xfanout1084 net1085 VGND VGND VPWR VPWR net1084 sky130_fd_sc_hd__clkbuf_2
Xfanout1095 _05428_ VGND VGND VPWR VPWR net1095 sky130_fd_sc_hd__buf_1
XFILLER_48_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05780_ _03249_ _03250_ _03260_ _03296_ VGND VGND VPWR VPWR _03297_ sky130_fd_sc_hd__or4_1
XFILLER_35_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13929_ clknet_leaf_73_clk _02558_ VGND VGND VPWR VPWR data_array.data1\[4\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07450_ net1222 _04685_ _04689_ net1173 VGND VGND VPWR VPWR _04691_ sky130_fd_sc_hd__a22o_1
XFILLER_179_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06401_ tag_array.tag0\[8\]\[19\] net1405 net1311 tag_array.tag0\[11\]\[19\] _03736_
+ VGND VGND VPWR VPWR _03737_ sky130_fd_sc_hd__a221o_1
X_07381_ data_array.data0\[1\]\[58\] net1545 net1449 data_array.data0\[2\]\[58\] VGND
+ VGND VPWR VPWR _04628_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_44_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09120_ net1063 net3506 net575 VGND VGND VPWR VPWR _00874_ sky130_fd_sc_hd__mux2_1
X_06332_ tag_array.tag0\[1\]\[13\] net1608 net1512 tag_array.tag0\[2\]\[13\] VGND
+ VGND VPWR VPWR _03674_ sky130_fd_sc_hd__a22o_1
XFILLER_163_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_844 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09051_ net1080 net2127 net416 VGND VGND VPWR VPWR _00805_ sky130_fd_sc_hd__mux2_1
X_06263_ _03610_ _03611_ VGND VGND VPWR VPWR _00152_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08002_ data_array.data1\[13\]\[51\] net1523 net1427 data_array.data1\[14\]\[51\]
+ VGND VGND VPWR VPWR _05192_ sky130_fd_sc_hd__a22o_1
XFILLER_117_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold501 data_array.data1\[9\]\[5\] VGND VGND VPWR VPWR net2152 sky130_fd_sc_hd__dlygate4sd3_1
X_06194_ tag_array.tag0\[0\]\[0\] net1404 net1310 tag_array.tag0\[3\]\[0\] _03548_
+ VGND VGND VPWR VPWR _03549_ sky130_fd_sc_hd__a221o_1
Xhold512 data_array.data1\[4\]\[51\] VGND VGND VPWR VPWR net2163 sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 data_array.data0\[4\]\[10\] VGND VGND VPWR VPWR net2174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 data_array.data0\[10\]\[5\] VGND VGND VPWR VPWR net2185 sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 tag_array.tag1\[1\]\[22\] VGND VGND VPWR VPWR net2196 sky130_fd_sc_hd__dlygate4sd3_1
Xhold556 tag_array.tag1\[1\]\[11\] VGND VGND VPWR VPWR net2207 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold567 data_array.data1\[2\]\[4\] VGND VGND VPWR VPWR net2218 sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 data_array.data1\[0\]\[47\] VGND VGND VPWR VPWR net2229 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09953_ net1018 net3459 net372 VGND VGND VPWR VPWR _01702_ sky130_fd_sc_hd__mux2_1
Xhold589 data_array.data0\[8\]\[24\] VGND VGND VPWR VPWR net2240 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_83_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08904_ net888 net4230 net435 VGND VGND VPWR VPWR _00661_ sky130_fd_sc_hd__mux2_1
XFILLER_44_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09884_ net933 net3555 net384 VGND VGND VPWR VPWR _01634_ sky130_fd_sc_hd__mux2_1
XFILLER_106_58 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1201 data_array.data1\[9\]\[59\] VGND VGND VPWR VPWR net2852 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1212 tag_array.tag0\[12\]\[14\] VGND VGND VPWR VPWR net2863 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_170_1075 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08835_ net2318 net904 net442 VGND VGND VPWR VPWR _00593_ sky130_fd_sc_hd__mux2_1
Xhold1223 data_array.data1\[12\]\[11\] VGND VGND VPWR VPWR net2874 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1234 tag_array.tag1\[12\]\[8\] VGND VGND VPWR VPWR net2885 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1245 data_array.data1\[3\]\[20\] VGND VGND VPWR VPWR net2896 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1256 data_array.data0\[6\]\[37\] VGND VGND VPWR VPWR net2907 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1267 data_array.data1\[11\]\[8\] VGND VGND VPWR VPWR net2918 sky130_fd_sc_hd__dlygate4sd3_1
X_08766_ net761 net2487 net452 VGND VGND VPWR VPWR _00525_ sky130_fd_sc_hd__mux2_1
Xhold1278 data_array.data0\[8\]\[21\] VGND VGND VPWR VPWR net2929 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05978_ data_array.rdata0\[49\] net850 net1147 VGND VGND VPWR VPWR _03446_ sky130_fd_sc_hd__o21a_1
Xhold1289 data_array.data1\[12\]\[10\] VGND VGND VPWR VPWR net2940 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07717_ data_array.data1\[12\]\[25\] net1331 net1237 data_array.data1\[15\]\[25\]
+ _04932_ VGND VGND VPWR VPWR _04933_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_140_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08697_ net2611 net734 net482 VGND VGND VPWR VPWR _00456_ sky130_fd_sc_hd__mux2_1
XFILLER_25_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07648_ net1176 _04865_ _04869_ net1224 VGND VGND VPWR VPWR _04871_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_101_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07579_ data_array.data1\[5\]\[12\] net1586 net1490 data_array.data1\[6\]\[12\] VGND
+ VGND VPWR VPWR _04808_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_24_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09318_ net707 net3013 net548 VGND VGND VPWR VPWR _01072_ sky130_fd_sc_hd__mux2_1
X_10590_ net1898 net1100 net468 VGND VGND VPWR VPWR _02335_ sky130_fd_sc_hd__mux2_1
XFILLER_21_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09249_ net782 net4020 net568 VGND VGND VPWR VPWR _01003_ sky130_fd_sc_hd__mux2_1
X_12260_ clknet_leaf_141_clk _01018_ VGND VGND VPWR VPWR tag_array.tag1\[14\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_147_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11211_ net931 net4073 net650 VGND VGND VPWR VPWR _02954_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12191_ clknet_leaf_159_clk _00999_ VGND VGND VPWR VPWR tag_array.tag0\[14\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_135_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11142_ net951 net4131 net551 VGND VGND VPWR VPWR _02885_ sky130_fd_sc_hd__mux2_1
XFILLER_107_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_164_3520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11073_ net1814 net971 net328 VGND VGND VPWR VPWR _02816_ sky130_fd_sc_hd__mux2_1
Xinput110 mem_rdata[1] VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_1
XFILLER_103_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput121 mem_rdata[2] VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_1
X_10024_ net990 net2928 net562 VGND VGND VPWR VPWR _01773_ sky130_fd_sc_hd__mux2_1
XFILLER_88_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput132 mem_rdata[3] VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_1
Xinput143 mem_rdata[4] VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_1
Xinput154 mem_rdata[5] VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_160_3439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2480 data_array.data1\[12\]\[40\] VGND VGND VPWR VPWR net4131 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2491 data_array.data0\[12\]\[52\] VGND VGND VPWR VPWR net4142 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1790 tag_array.tag0\[7\]\[21\] VGND VGND VPWR VPWR net3441 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_147_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11975_ clknet_leaf_61_clk _00783_ VGND VGND VPWR VPWR data_array.data0\[4\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
X_13714_ clknet_leaf_117_clk _02343_ VGND VGND VPWR VPWR data_array.data1\[1\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_10926_ net1038 net4338 net531 VGND VGND VPWR VPWR _02671_ sky130_fd_sc_hd__mux2_1
XFILLER_71_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13645_ clknet_leaf_197_clk _02274_ VGND VGND VPWR VPWR data_array.data1\[15\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_10857_ net1056 net3817 net516 VGND VGND VPWR VPWR _02602_ sky130_fd_sc_hd__mux2_1
XFILLER_31_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13576_ clknet_leaf_5_clk _02205_ VGND VGND VPWR VPWR data_array.data0\[9\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10788_ net2212 net1079 net503 VGND VGND VPWR VPWR _02533_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12527_ clknet_leaf_141_clk _01221_ VGND VGND VPWR VPWR tag_array.tag1\[11\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_858 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12458_ clknet_leaf_118_clk _01152_ VGND VGND VPWR VPWR data_array.data1\[9\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_10_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11409_ clknet_leaf_129_clk _00219_ VGND VGND VPWR VPWR tag_array.tag1\[7\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_160_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12389_ clknet_leaf_104_clk _01083_ VGND VGND VPWR VPWR data_array.data0\[14\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_184_3907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_184_3918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14128_ clknet_leaf_109_clk _02757_ VGND VGND VPWR VPWR data_array.data0\[1\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_98_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06950_ data_array.data0\[9\]\[19\] net1582 net1486 data_array.data0\[10\]\[19\]
+ VGND VGND VPWR VPWR _04236_ sky130_fd_sc_hd__a22o_1
X_14059_ clknet_leaf_256_clk _02688_ VGND VGND VPWR VPWR data_array.data1\[6\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_67_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05901_ data_array.rdata1\[23\] net830 net840 VGND VGND VPWR VPWR _03395_ sky130_fd_sc_hd__a21o_1
XFILLER_140_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06881_ data_array.data0\[12\]\[13\] net1361 net1267 data_array.data0\[15\]\[13\]
+ _04172_ VGND VGND VPWR VPWR _04173_ sky130_fd_sc_hd__a221o_1
X_08620_ net743 net3700 net525 VGND VGND VPWR VPWR _00379_ sky130_fd_sc_hd__mux2_1
X_05832_ _03348_ data_array.rdata0\[0\] net827 VGND VGND VPWR VPWR _03349_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_85_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08551_ net751 net3216 net589 VGND VGND VPWR VPWR _00319_ sky130_fd_sc_hd__mux2_1
X_05763_ fsm.tag_out1\[23\] net24 VGND VGND VPWR VPWR _03280_ sky130_fd_sc_hd__and2b_1
XFILLER_36_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07502_ data_array.data1\[5\]\[5\] net1551 net1455 data_array.data1\[6\]\[5\] VGND
+ VGND VPWR VPWR _04738_ sky130_fd_sc_hd__a22o_1
XFILLER_74_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08482_ net1564 net1200 VGND VGND VPWR VPWR _05558_ sky130_fd_sc_hd__nand2_1
XFILLER_50_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05694_ _03207_ _03208_ _03209_ _03210_ VGND VGND VPWR VPWR _03211_ sky130_fd_sc_hd__or4_4
X_07433_ data_array.data0\[4\]\[63\] net1366 net1272 data_array.data0\[7\]\[63\] _04674_
+ VGND VGND VPWR VPWR _04675_ sky130_fd_sc_hd__a221o_1
XFILLER_50_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_77_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07364_ data_array.data0\[13\]\[57\] net1541 net1445 data_array.data0\[14\]\[57\]
+ VGND VGND VPWR VPWR _04612_ sky130_fd_sc_hd__a22o_1
XFILLER_22_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09103_ net872 net3867 net414 VGND VGND VPWR VPWR _00857_ sky130_fd_sc_hd__mux2_1
X_06315_ tag_array.tag0\[4\]\[11\] net1402 net1308 tag_array.tag0\[7\]\[11\] _03658_
+ VGND VGND VPWR VPWR _03659_ sky130_fd_sc_hd__a221o_1
XFILLER_148_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07295_ net1619 _04543_ _04547_ net1193 VGND VGND VPWR VPWR _04550_ sky130_fd_sc_hd__a22o_1
XFILLER_136_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09034_ net2063 net888 net419 VGND VGND VPWR VPWR _00789_ sky130_fd_sc_hd__mux2_1
X_06246_ tag_array.tag0\[9\]\[5\] net1608 net1512 tag_array.tag0\[10\]\[5\] VGND VGND
+ VPWR VPWR _03596_ sky130_fd_sc_hd__a22o_1
XFILLER_163_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold320 data_array.data1\[8\]\[34\] VGND VGND VPWR VPWR net1971 sky130_fd_sc_hd__dlygate4sd3_1
Xhold331 data_array.data1\[8\]\[10\] VGND VGND VPWR VPWR net1982 sky130_fd_sc_hd__dlygate4sd3_1
X_06177_ tag_array.valid1\[12\] net1369 net1275 tag_array.valid1\[15\] _03532_ VGND
+ VGND VPWR VPWR _03533_ sky130_fd_sc_hd__a221o_1
XFILLER_116_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold342 data_array.data1\[1\]\[49\] VGND VGND VPWR VPWR net1993 sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 data_array.data1\[2\]\[36\] VGND VGND VPWR VPWR net2004 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold364 tag_array.tag1\[1\]\[6\] VGND VGND VPWR VPWR net2015 sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 data_array.data0\[4\]\[1\] VGND VGND VPWR VPWR net2026 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_57_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold386 data_array.data1\[1\]\[20\] VGND VGND VPWR VPWR net2037 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout800 net803 VGND VGND VPWR VPWR net800 sky130_fd_sc_hd__buf_4
XFILLER_120_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold397 data_array.data0\[1\]\[16\] VGND VGND VPWR VPWR net2048 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout811 net815 VGND VGND VPWR VPWR net811 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_86_Right_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09936_ net1084 net4025 net370 VGND VGND VPWR VPWR _01685_ sky130_fd_sc_hd__mux2_1
Xfanout822 net823 VGND VGND VPWR VPWR net822 sky130_fd_sc_hd__buf_1
Xfanout833 net834 VGND VGND VPWR VPWR net833 sky130_fd_sc_hd__buf_8
Xfanout844 net845 VGND VGND VPWR VPWR net844 sky130_fd_sc_hd__buf_8
Xfanout855 _05554_ VGND VGND VPWR VPWR net855 sky130_fd_sc_hd__clkbuf_2
Xfanout866 _05542_ VGND VGND VPWR VPWR net866 sky130_fd_sc_hd__clkbuf_2
XFILLER_58_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_142_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout877 _05536_ VGND VGND VPWR VPWR net877 sky130_fd_sc_hd__dlymetal6s2s_1
X_09867_ net1002 net4502 net381 VGND VGND VPWR VPWR _01617_ sky130_fd_sc_hd__mux2_1
XFILLER_85_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1020 data_array.data0\[0\]\[39\] VGND VGND VPWR VPWR net2671 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout888 _05530_ VGND VGND VPWR VPWR net888 sky130_fd_sc_hd__clkbuf_2
Xfanout899 _05526_ VGND VGND VPWR VPWR net899 sky130_fd_sc_hd__buf_1
Xhold1031 data_array.data0\[9\]\[8\] VGND VGND VPWR VPWR net2682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1042 data_array.data1\[15\]\[7\] VGND VGND VPWR VPWR net2693 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08818_ net2626 net973 net442 VGND VGND VPWR VPWR _00576_ sky130_fd_sc_hd__mux2_1
XFILLER_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1053 tag_array.tag1\[12\]\[15\] VGND VGND VPWR VPWR net2704 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1064 data_array.data0\[5\]\[58\] VGND VGND VPWR VPWR net2715 sky130_fd_sc_hd__dlygate4sd3_1
X_09798_ net1018 net4573 net388 VGND VGND VPWR VPWR _01549_ sky130_fd_sc_hd__mux2_1
XFILLER_93_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1075 tag_array.tag0\[13\]\[11\] VGND VGND VPWR VPWR net2726 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1086 data_array.data0\[12\]\[61\] VGND VGND VPWR VPWR net2737 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1097 tag_array.tag1\[2\]\[0\] VGND VGND VPWR VPWR net2748 sky130_fd_sc_hd__dlygate4sd3_1
X_08749_ net729 net2674 net463 VGND VGND VPWR VPWR _00508_ sky130_fd_sc_hd__mux2_1
XFILLER_27_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_5_23__f_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_5_23__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_73_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11760_ clknet_leaf_240_clk _00568_ VGND VGND VPWR VPWR data_array.data0\[8\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_158_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_95_Right_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10711_ net2587 net875 net483 VGND VGND VPWR VPWR _02456_ sky130_fd_sc_hd__mux2_1
X_11691_ clknet_leaf_133_clk _00499_ VGND VGND VPWR VPWR tag_array.tag1\[15\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10642_ net2628 net892 net469 VGND VGND VPWR VPWR _02387_ sky130_fd_sc_hd__mux2_1
X_13430_ clknet_leaf_242_clk _02060_ VGND VGND VPWR VPWR data_array.data1\[8\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_157_3390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13361_ clknet_leaf_179_clk _01991_ VGND VGND VPWR VPWR tag_array.tag0\[2\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_139_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_118_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10573_ net915 net3311 net461 VGND VGND VPWR VPWR _02318_ sky130_fd_sc_hd__mux2_1
XFILLER_166_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12312_ clknet_leaf_103_clk _01070_ VGND VGND VPWR VPWR tag_array.tag1\[12\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_13292_ clknet_leaf_5_clk _01922_ VGND VGND VPWR VPWR data_array.data0\[10\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_846 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12243_ clknet_leaf_96_clk _01001_ VGND VGND VPWR VPWR tag_array.tag1\[14\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_114_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12174_ clknet_leaf_154_clk _00982_ VGND VGND VPWR VPWR tag_array.tag0\[14\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_131_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11125_ net1016 net2890 net545 VGND VGND VPWR VPWR _02868_ sky130_fd_sc_hd__mux2_1
XFILLER_77_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11056_ net2725 net1036 net329 VGND VGND VPWR VPWR _02799_ sky130_fd_sc_hd__mux2_1
X_10007_ net1057 net2858 net558 VGND VGND VPWR VPWR _01756_ sky130_fd_sc_hd__mux2_1
XFILLER_3_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11958_ clknet_leaf_264_clk _00766_ VGND VGND VPWR VPWR data_array.data0\[4\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_83_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_177_3755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_177_3766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10909_ net1104 net4410 net526 VGND VGND VPWR VPWR _02654_ sky130_fd_sc_hd__mux2_1
XFILLER_60_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11889_ clknet_leaf_238_clk _00697_ VGND VGND VPWR VPWR data_array.data0\[5\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_73_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13628_ clknet_leaf_10_clk _02257_ VGND VGND VPWR VPWR data_array.data0\[9\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_15_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13559_ clknet_leaf_9_clk _02188_ VGND VGND VPWR VPWR data_array.data1\[0\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06100_ data_array.rdata0\[15\] net1139 net1114 data_array.rdata1\[15\] VGND VGND
+ VPWR VPWR net269 sky130_fd_sc_hd__a22o_1
XFILLER_8_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07080_ data_array.data0\[5\]\[31\] net1574 net1478 data_array.data0\[6\]\[31\] VGND
+ VGND VPWR VPWR _04354_ sky130_fd_sc_hd__a22o_1
XFILLER_172_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06031_ net1160 net1137 net1118 net26 VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__o31a_1
XFILLER_161_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_327 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_262_clk clknet_5_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_262_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_99_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07982_ data_array.data1\[1\]\[49\] net1572 net1476 data_array.data1\[2\]\[49\] VGND
+ VGND VPWR VPWR _05174_ sky130_fd_sc_hd__a22o_1
XFILLER_99_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06933_ net1214 _04215_ _04219_ net1166 VGND VGND VPWR VPWR _04221_ sky130_fd_sc_hd__a22o_1
X_09721_ net704 net3513 net611 VGND VGND VPWR VPWR _01473_ sky130_fd_sc_hd__mux2_1
XFILLER_68_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_52_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09652_ net781 net3714 net612 VGND VGND VPWR VPWR _01404_ sky130_fd_sc_hd__mux2_1
X_06864_ data_array.data0\[5\]\[11\] net1568 net1472 data_array.data0\[6\]\[11\] VGND
+ VGND VPWR VPWR _04158_ sky130_fd_sc_hd__a22o_1
XFILLER_82_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08603_ net710 net4613 net527 VGND VGND VPWR VPWR _00362_ sky130_fd_sc_hd__mux2_1
X_05815_ _03328_ _03329_ _03330_ _03331_ VGND VGND VPWR VPWR _03332_ sky130_fd_sc_hd__or4_1
X_09583_ net1019 net4058 net397 VGND VGND VPWR VPWR _01335_ sky130_fd_sc_hd__mux2_1
X_06795_ data_array.data0\[0\]\[5\] net1360 net1266 data_array.data0\[3\]\[5\] _04094_
+ VGND VGND VPWR VPWR _04095_ sky130_fd_sc_hd__a221o_1
X_08534_ net1559 net1200 net814 net1707 VGND VGND VPWR VPWR _00306_ sky130_fd_sc_hd__a31o_1
X_05746_ fsm.tag_out1\[21\] net21 VGND VGND VPWR VPWR _03263_ sky130_fd_sc_hd__and2b_1
XFILLER_35_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08465_ net2496 net856 net688 VGND VGND VPWR VPWR _00284_ sky130_fd_sc_hd__mux2_1
X_05677_ fsm.tag_out0\[9\] net8 VGND VGND VPWR VPWR _03194_ sky130_fd_sc_hd__and2b_1
XFILLER_24_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07416_ net1196 _04653_ _04657_ net1622 VGND VGND VPWR VPWR _04660_ sky130_fd_sc_hd__a22o_1
XFILLER_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08396_ net2146 net948 net693 VGND VGND VPWR VPWR _00261_ sky130_fd_sc_hd__mux2_1
XFILLER_10_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07347_ data_array.data0\[8\]\[55\] net1343 net1249 data_array.data0\[11\]\[55\]
+ _04596_ VGND VGND VPWR VPWR _04597_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_98_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07278_ data_array.data0\[1\]\[49\] net1571 net1475 data_array.data0\[2\]\[49\] VGND
+ VGND VPWR VPWR _04534_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_59_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09017_ net2924 net956 net422 VGND VGND VPWR VPWR _00772_ sky130_fd_sc_hd__mux2_1
XFILLER_128_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06229_ net1221 _03575_ _03579_ net1172 VGND VGND VPWR VPWR _03581_ sky130_fd_sc_hd__a22o_1
XFILLER_163_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold150 tag_array.tag1\[0\]\[16\] VGND VGND VPWR VPWR net1801 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold161 tag_array.tag1\[1\]\[5\] VGND VGND VPWR VPWR net1812 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 data_array.data1\[0\]\[4\] VGND VGND VPWR VPWR net1823 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 data_array.data0\[0\]\[47\] VGND VGND VPWR VPWR net1834 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_253_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_253_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold194 tag_array.tag1\[0\]\[2\] VGND VGND VPWR VPWR net1845 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout1606 net1612 VGND VGND VPWR VPWR net1606 sky130_fd_sc_hd__buf_2
Xfanout1617 net1627 VGND VGND VPWR VPWR net1617 sky130_fd_sc_hd__buf_2
Xfanout630 net632 VGND VGND VPWR VPWR net630 sky130_fd_sc_hd__buf_4
XFILLER_104_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1628 net1629 VGND VGND VPWR VPWR net1628 sky130_fd_sc_hd__clkbuf_4
Xfanout641 net644 VGND VGND VPWR VPWR net641 sky130_fd_sc_hd__clkbuf_4
Xfanout1639 net1642 VGND VGND VPWR VPWR net1639 sky130_fd_sc_hd__clkbuf_8
Xfanout652 net654 VGND VGND VPWR VPWR net652 sky130_fd_sc_hd__clkbuf_8
X_09919_ net732 net2683 net603 VGND VGND VPWR VPWR _01669_ sky130_fd_sc_hd__mux2_1
Xfanout663 net666 VGND VGND VPWR VPWR net663 sky130_fd_sc_hd__clkbuf_8
Xfanout674 net676 VGND VGND VPWR VPWR net674 sky130_fd_sc_hd__clkbuf_4
Xfanout685 _05548_ VGND VGND VPWR VPWR net685 sky130_fd_sc_hd__buf_4
X_12930_ clknet_leaf_10_clk _01624_ VGND VGND VPWR VPWR data_array.data0\[13\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout696 net697 VGND VGND VPWR VPWR net696 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_124_Left_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12861_ clknet_leaf_55_clk _01555_ VGND VGND VPWR VPWR data_array.data0\[12\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_160_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11812_ clknet_leaf_50_clk _00620_ VGND VGND VPWR VPWR data_array.data0\[7\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12792_ clknet_leaf_104_clk _01486_ VGND VGND VPWR VPWR tag_array.tag1\[10\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11743_ clknet_leaf_60_clk _00551_ VGND VGND VPWR VPWR data_array.data0\[8\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_155_3338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_155_3349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14462_ clknet_leaf_261_clk _03085_ VGND VGND VPWR VPWR data_array.data1\[7\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11674_ clknet_leaf_98_clk _00482_ VGND VGND VPWR VPWR tag_array.tag1\[1\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_12_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13413_ clknet_leaf_76_clk _02043_ VGND VGND VPWR VPWR data_array.data1\[8\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_172_3663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10625_ net2997 net960 net469 VGND VGND VPWR VPWR _02370_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_172_3674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14393_ clknet_leaf_43_clk _03016_ VGND VGND VPWR VPWR data_array.data1\[10\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_133_Left_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10556_ net981 net4026 net453 VGND VGND VPWR VPWR _02301_ sky130_fd_sc_hd__mux2_1
X_13344_ clknet_leaf_11_clk _01974_ VGND VGND VPWR VPWR data_array.data0\[10\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_133_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10487_ net998 net4499 net345 VGND VGND VPWR VPWR _02232_ sky130_fd_sc_hd__mux2_1
X_13275_ clknet_leaf_90_clk _01905_ VGND VGND VPWR VPWR data_array.data0\[11\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_142_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12226_ clknet_leaf_148_clk _00179_ VGND VGND VPWR VPWR fsm.tag_out1\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_184_Right_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_244_clk clknet_5_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_244_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12157_ clknet_leaf_173_clk _00965_ VGND VGND VPWR VPWR tag_array.tag0\[13\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_151_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11108_ net1086 net3979 net541 VGND VGND VPWR VPWR _02851_ sky130_fd_sc_hd__mux2_1
XFILLER_68_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12088_ clknet_leaf_8_clk _00896_ VGND VGND VPWR VPWR data_array.data1\[14\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_96_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_142_Left_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11039_ net3997 net1105 net328 VGND VGND VPWR VPWR _02782_ sky130_fd_sc_hd__mux2_1
XFILLER_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_179_3806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_536 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06580_ net1207 _03893_ _03897_ net1633 VGND VGND VPWR VPWR _03900_ sky130_fd_sc_hd__a22o_1
XFILLER_18_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08250_ net719 net2233 net799 VGND VGND VPWR VPWR _00214_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_151_Left_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07201_ data_array.data0\[5\]\[42\] net1579 net1483 data_array.data0\[6\]\[42\] VGND
+ VGND VPWR VPWR _04464_ sky130_fd_sc_hd__a22o_1
X_08181_ _03511_ _03519_ VGND VGND VPWR VPWR _05352_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_31_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07132_ _04400_ _04401_ VGND VGND VPWR VPWR _00028_ sky130_fd_sc_hd__or2_1
XFILLER_173_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07063_ data_array.data0\[4\]\[29\] net1380 net1286 data_array.data0\[7\]\[29\] _04338_
+ VGND VGND VPWR VPWR _04339_ sky130_fd_sc_hd__a221o_1
XFILLER_161_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput200 net200 VGND VGND VPWR VPWR cpu_rdata[41] sky130_fd_sc_hd__buf_2
Xoutput211 net211 VGND VGND VPWR VPWR cpu_rdata[51] sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_93_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06014_ data_array.rdata0\[61\] net849 net1145 VGND VGND VPWR VPWR _03470_ sky130_fd_sc_hd__o21a_1
Xoutput222 net222 VGND VGND VPWR VPWR cpu_rdata[61] sky130_fd_sc_hd__buf_2
Xoutput233 net233 VGND VGND VPWR VPWR mem_addr[12] sky130_fd_sc_hd__buf_2
Xoutput244 net244 VGND VGND VPWR VPWR mem_addr[22] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput255 net255 VGND VGND VPWR VPWR mem_addr[3] sky130_fd_sc_hd__buf_2
Xoutput266 net266 VGND VGND VPWR VPWR mem_wdata[12] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_151_Right_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_235_clk clknet_5_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_235_clk
+ sky130_fd_sc_hd__clkbuf_8
Xoutput277 net277 VGND VGND VPWR VPWR mem_wdata[22] sky130_fd_sc_hd__buf_2
Xoutput288 net288 VGND VGND VPWR VPWR mem_wdata[32] sky130_fd_sc_hd__buf_2
Xoutput299 net299 VGND VGND VPWR VPWR mem_wdata[42] sky130_fd_sc_hd__buf_2
XFILLER_99_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_160_Left_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07965_ data_array.data1\[0\]\[47\] net1397 net1303 data_array.data1\[3\]\[47\] _05158_
+ VGND VGND VPWR VPWR _05159_ sky130_fd_sc_hd__a221o_1
XFILLER_74_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09704_ net770 net4149 net610 VGND VGND VPWR VPWR _01456_ sky130_fd_sc_hd__mux2_1
X_06916_ data_array.data0\[4\]\[16\] net1356 net1262 data_array.data0\[7\]\[16\] _04204_
+ VGND VGND VPWR VPWR _04205_ sky130_fd_sc_hd__a221o_1
XFILLER_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07896_ data_array.data1\[13\]\[41\] net1525 net1429 data_array.data1\[14\]\[41\]
+ VGND VGND VPWR VPWR _05096_ sky130_fd_sc_hd__a22o_1
XFILLER_110_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09635_ net748 net3961 net616 VGND VGND VPWR VPWR _01387_ sky130_fd_sc_hd__mux2_1
XFILLER_56_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06847_ data_array.data0\[9\]\[10\] net1601 net1505 data_array.data0\[10\]\[10\]
+ VGND VGND VPWR VPWR _04142_ sky130_fd_sc_hd__a22o_1
XFILLER_71_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09566_ net1085 net3444 net394 VGND VGND VPWR VPWR _01318_ sky130_fd_sc_hd__mux2_1
X_06778_ net1202 _04073_ _04077_ net1628 VGND VGND VPWR VPWR _04080_ sky130_fd_sc_hd__a22o_1
X_05729_ net2 fsm.tag_out1\[3\] VGND VGND VPWR VPWR _03246_ sky130_fd_sc_hd__xor2_1
X_08517_ net1716 net604 VGND VGND VPWR VPWR _00300_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_137_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09497_ net738 net2393 net626 VGND VGND VPWR VPWR _01250_ sky130_fd_sc_hd__mux2_1
XFILLER_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08448_ net152 net87 net1643 VGND VGND VPWR VPWR _05535_ sky130_fd_sc_hd__mux2_1
XFILLER_11_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1050 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08379_ net127 net62 net1639 VGND VGND VPWR VPWR _05489_ sky130_fd_sc_hd__mux2_1
XFILLER_109_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10410_ net1976 net1015 net670 VGND VGND VPWR VPWR _02156_ sky130_fd_sc_hd__mux2_1
XFILLER_139_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11390_ clknet_leaf_194_clk _00200_ VGND VGND VPWR VPWR tag_array.tag1\[7\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_109_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_150_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10341_ net735 net4100 net591 VGND VGND VPWR VPWR _02088_ sky130_fd_sc_hd__mux2_1
XFILLER_87_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13060_ clknet_leaf_35_clk _01754_ VGND VGND VPWR VPWR data_array.data1\[13\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_105_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10272_ net1852 net1075 net640 VGND VGND VPWR VPWR _02019_ sky130_fd_sc_hd__mux2_1
XFILLER_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12011_ clknet_leaf_228_clk _00819_ VGND VGND VPWR VPWR data_array.data0\[6\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_105_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_226_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_226_clk
+ sky130_fd_sc_hd__clkbuf_8
Xfanout1403 net1406 VGND VGND VPWR VPWR net1403 sky130_fd_sc_hd__clkbuf_4
Xfanout1414 net1416 VGND VGND VPWR VPWR net1414 sky130_fd_sc_hd__clkbuf_4
Xfanout1425 net1447 VGND VGND VPWR VPWR net1425 sky130_fd_sc_hd__clkbuf_2
XFILLER_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1436 net1437 VGND VGND VPWR VPWR net1436 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1447 net1518 VGND VGND VPWR VPWR net1447 sky130_fd_sc_hd__clkbuf_4
Xfanout1458 net1518 VGND VGND VPWR VPWR net1458 sky130_fd_sc_hd__buf_2
Xfanout460 net465 VGND VGND VPWR VPWR net460 sky130_fd_sc_hd__buf_4
Xfanout1469 net1470 VGND VGND VPWR VPWR net1469 sky130_fd_sc_hd__clkbuf_2
Xfanout471 net474 VGND VGND VPWR VPWR net471 sky130_fd_sc_hd__clkbuf_8
Xfanout482 net489 VGND VGND VPWR VPWR net482 sky130_fd_sc_hd__buf_6
X_13962_ clknet_leaf_251_clk _02591_ VGND VGND VPWR VPWR data_array.data1\[5\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout493 net494 VGND VGND VPWR VPWR net493 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_109_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12913_ clknet_leaf_246_clk _01607_ VGND VGND VPWR VPWR data_array.data0\[13\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13893_ clknet_leaf_211_clk _02522_ VGND VGND VPWR VPWR data_array.data1\[3\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_126_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12844_ clknet_leaf_104_clk _01538_ VGND VGND VPWR VPWR data_array.data0\[12\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_17_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ clknet_leaf_153_clk _01469_ VGND VGND VPWR VPWR tag_array.tag0\[6\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_11726_ clknet_leaf_108_clk _00534_ VGND VGND VPWR VPWR tag_array.tag0\[9\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14445_ clknet_leaf_39_clk _03068_ VGND VGND VPWR VPWR data_array.data1\[7\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_11657_ clknet_leaf_128_clk _00465_ VGND VGND VPWR VPWR tag_array.tag1\[2\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_174_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10608_ net2037 net1030 net475 VGND VGND VPWR VPWR _02353_ sky130_fd_sc_hd__mux2_1
XFILLER_11_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14376_ clknet_leaf_259_clk _02999_ VGND VGND VPWR VPWR data_array.data1\[10\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_11588_ clknet_leaf_194_clk _00396_ VGND VGND VPWR VPWR tag_array.tag1\[4\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold908 data_array.data1\[13\]\[62\] VGND VGND VPWR VPWR net2559 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_923 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13327_ clknet_leaf_116_clk _01957_ VGND VGND VPWR VPWR data_array.data0\[10\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_182_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10539_ net1050 net3401 net461 VGND VGND VPWR VPWR _02284_ sky130_fd_sc_hd__mux2_1
Xhold919 tag_array.tag0\[14\]\[6\] VGND VGND VPWR VPWR net2570 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_109_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13258_ clknet_leaf_38_clk _01888_ VGND VGND VPWR VPWR data_array.data0\[11\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_171_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_217_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_217_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12209_ clknet_leaf_148_clk _00138_ VGND VGND VPWR VPWR fsm.tag_out0\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_1026 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13189_ clknet_leaf_254_clk _00082_ VGND VGND VPWR VPWR data_array.rdata1\[26\] sky130_fd_sc_hd__dfxtp_1
Xhold2309 data_array.data1\[10\]\[50\] VGND VGND VPWR VPWR net3960 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1608 data_array.data0\[12\]\[50\] VGND VGND VPWR VPWR net3259 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1619 data_array.data0\[4\]\[39\] VGND VGND VPWR VPWR net3270 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07750_ data_array.data1\[8\]\[28\] net1349 net1255 data_array.data1\[11\]\[28\]
+ _04962_ VGND VGND VPWR VPWR _04963_ sky130_fd_sc_hd__a221o_1
XFILLER_49_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06701_ net1633 _04003_ _04007_ net1207 VGND VGND VPWR VPWR _04010_ sky130_fd_sc_hd__a22o_1
XFILLER_38_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07681_ net1222 _04895_ _04899_ net1173 VGND VGND VPWR VPWR _04901_ sky130_fd_sc_hd__a22o_1
XFILLER_53_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06632_ tag_array.tag1\[12\]\[15\] net1403 net1309 tag_array.tag1\[15\]\[15\] _03946_
+ VGND VGND VPWR VPWR _03947_ sky130_fd_sc_hd__a221o_1
X_09420_ net985 net3542 net585 VGND VGND VPWR VPWR _01173_ sky130_fd_sc_hd__mux2_1
XFILLER_53_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09351_ net998 net3984 net406 VGND VGND VPWR VPWR _01104_ sky130_fd_sc_hd__mux2_1
X_06563_ tag_array.tag1\[5\]\[9\] net1607 net1511 tag_array.tag1\[6\]\[9\] VGND VGND
+ VPWR VPWR _03884_ sky130_fd_sc_hd__a22o_1
XFILLER_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08302_ net1127 _05437_ VGND VGND VPWR VPWR _05438_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_47_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09282_ net751 net3648 net565 VGND VGND VPWR VPWR _01036_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06494_ _03820_ _03821_ VGND VGND VPWR VPWR _00173_ sky130_fd_sc_hd__or2_2
XFILLER_139_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08233_ net1650 net1163 net13 VGND VGND VPWR VPWR _05390_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_95_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08164_ net1207 _05333_ _05337_ net1633 VGND VGND VPWR VPWR _05340_ sky130_fd_sc_hd__a22o_1
XFILLER_162_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07115_ data_array.data0\[9\]\[34\] net1531 net1435 data_array.data0\[10\]\[34\]
+ VGND VGND VPWR VPWR _04386_ sky130_fd_sc_hd__a22o_1
X_08095_ data_array.data1\[12\]\[59\] net1381 net1287 data_array.data1\[15\]\[59\]
+ _05276_ VGND VGND VPWR VPWR _05277_ sky130_fd_sc_hd__a221o_1
XFILLER_134_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload70 clknet_leaf_236_clk VGND VGND VPWR VPWR clkload70/Y sky130_fd_sc_hd__inv_12
XFILLER_161_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07046_ data_array.data0\[8\]\[28\] net1351 net1257 data_array.data0\[11\]\[28\]
+ _04322_ VGND VGND VPWR VPWR _04323_ sky130_fd_sc_hd__a221o_1
Xclkload81 clknet_leaf_40_clk VGND VGND VPWR VPWR clkload81/Y sky130_fd_sc_hd__bufinv_16
Xclkload92 clknet_leaf_65_clk VGND VGND VPWR VPWR clkload92/Y sky130_fd_sc_hd__clkinv_8
XFILLER_161_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_208_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_208_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_88_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2810 tag_array.tag1\[4\]\[9\] VGND VGND VPWR VPWR net4461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2821 data_array.data0\[14\]\[47\] VGND VGND VPWR VPWR net4472 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_125_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2832 data_array.data0\[5\]\[32\] VGND VGND VPWR VPWR net4483 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_778 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08997_ net2138 net1036 net423 VGND VGND VPWR VPWR _00752_ sky130_fd_sc_hd__mux2_1
Xhold2843 data_array.data1\[15\]\[3\] VGND VGND VPWR VPWR net4494 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2854 data_array.data1\[7\]\[38\] VGND VGND VPWR VPWR net4505 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2865 tag_array.tag1\[6\]\[7\] VGND VGND VPWR VPWR net4516 sky130_fd_sc_hd__dlygate4sd3_1
X_07948_ data_array.data1\[8\]\[46\] net1337 net1243 data_array.data1\[11\]\[46\]
+ _05142_ VGND VGND VPWR VPWR _05143_ sky130_fd_sc_hd__a221o_1
Xhold2876 tag_array.tag0\[7\]\[24\] VGND VGND VPWR VPWR net4527 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2887 data_array.data1\[10\]\[22\] VGND VGND VPWR VPWR net4538 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2898 data_array.data1\[15\]\[1\] VGND VGND VPWR VPWR net4549 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07879_ net1217 _05075_ _05079_ net1169 VGND VGND VPWR VPWR _05081_ sky130_fd_sc_hd__a22o_1
XFILLER_71_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09618_ net877 net3174 net397 VGND VGND VPWR VPWR _01370_ sky130_fd_sc_hd__mux2_1
X_10890_ net925 net3674 net514 VGND VGND VPWR VPWR _02635_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_104_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09549_ net732 net3544 net618 VGND VGND VPWR VPWR _01302_ sky130_fd_sc_hd__mux2_1
XFILLER_12_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12560_ clknet_leaf_108_clk _01254_ VGND VGND VPWR VPWR tag_array.tag0\[11\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_157_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11511_ clknet_leaf_104_clk _00319_ VGND VGND VPWR VPWR tag_array.tag1\[9\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_169_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12491_ clknet_leaf_43_clk _01185_ VGND VGND VPWR VPWR data_array.data1\[9\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_141_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14230_ clknet_leaf_41_clk _02859_ VGND VGND VPWR VPWR data_array.data1\[12\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_156_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11442_ clknet_leaf_34_clk _00252_ VGND VGND VPWR VPWR data_array.data0\[0\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_172_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11373_ net1647 net3765 net628 VGND VGND VPWR VPWR _03116_ sky130_fd_sc_hd__mux2_1
X_14161_ clknet_leaf_62_clk _02790_ VGND VGND VPWR VPWR data_array.data0\[2\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_166_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10324_ net2073 net864 net637 VGND VGND VPWR VPWR _02071_ sky130_fd_sc_hd__mux2_1
X_13112_ clknet_leaf_192_clk _01806_ VGND VGND VPWR VPWR data_array.data1\[13\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14092_ clknet_leaf_71_clk _02721_ VGND VGND VPWR VPWR data_array.data0\[1\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13043_ clknet_leaf_207_clk _01737_ VGND VGND VPWR VPWR data_array.data0\[3\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
X_10255_ net722 net2646 net596 VGND VGND VPWR VPWR _02002_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_167_3562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_3573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1200 net1201 VGND VGND VPWR VPWR net1200 sky130_fd_sc_hd__buf_4
XFILLER_59_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1211 net1212 VGND VGND VPWR VPWR net1211 sky130_fd_sc_hd__buf_4
XFILLER_105_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1222 net1223 VGND VGND VPWR VPWR net1222 sky130_fd_sc_hd__buf_4
X_10186_ net1061 net3422 net360 VGND VGND VPWR VPWR _01933_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1233 net1234 VGND VGND VPWR VPWR net1233 sky130_fd_sc_hd__buf_4
XFILLER_182_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1244 net1245 VGND VGND VPWR VPWR net1244 sky130_fd_sc_hd__clkbuf_4
XFILLER_79_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1255 net1257 VGND VGND VPWR VPWR net1255 sky130_fd_sc_hd__clkbuf_4
XFILLER_121_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1266 net1270 VGND VGND VPWR VPWR net1266 sky130_fd_sc_hd__clkbuf_4
Xfanout1277 net1281 VGND VGND VPWR VPWR net1277 sky130_fd_sc_hd__clkbuf_4
Xfanout1288 net1289 VGND VGND VPWR VPWR net1288 sky130_fd_sc_hd__clkbuf_2
Xfanout1299 net1300 VGND VGND VPWR VPWR net1299 sky130_fd_sc_hd__clkbuf_4
XFILLER_19_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13945_ clknet_leaf_55_clk _02574_ VGND VGND VPWR VPWR data_array.data1\[4\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_93_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_995 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13876_ clknet_leaf_83_clk _02505_ VGND VGND VPWR VPWR data_array.data1\[3\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12827_ clknet_leaf_232_clk _01521_ VGND VGND VPWR VPWR tag_array.tag1\[0\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12758_ clknet_leaf_166_clk _01452_ VGND VGND VPWR VPWR tag_array.tag0\[6\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11709_ clknet_leaf_106_clk _00517_ VGND VGND VPWR VPWR tag_array.tag0\[9\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_12689_ clknet_leaf_144_clk _01383_ VGND VGND VPWR VPWR tag_array.tag0\[8\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14428_ clknet_leaf_86_clk _03051_ VGND VGND VPWR VPWR data_array.data1\[7\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_156_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold705 tag_array.tag1\[12\]\[18\] VGND VGND VPWR VPWR net2356 sky130_fd_sc_hd__dlygate4sd3_1
X_14359_ clknet_leaf_58_clk _02982_ VGND VGND VPWR VPWR data_array.data1\[10\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold716 tag_array.tag1\[3\]\[8\] VGND VGND VPWR VPWR net2367 sky130_fd_sc_hd__dlygate4sd3_1
Xhold727 data_array.data0\[12\]\[15\] VGND VGND VPWR VPWR net2378 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_956 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold738 tag_array.tag1\[5\]\[22\] VGND VGND VPWR VPWR net2389 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold749 data_array.data0\[12\]\[60\] VGND VGND VPWR VPWR net2400 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08920_ net1085 net2966 net426 VGND VGND VPWR VPWR _00676_ sky130_fd_sc_hd__mux2_1
Xhold2106 tag_array.tag1\[12\]\[23\] VGND VGND VPWR VPWR net3757 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2117 tag_array.tag1\[6\]\[24\] VGND VGND VPWR VPWR net3768 sky130_fd_sc_hd__dlygate4sd3_1
X_08851_ net1102 net2334 net436 VGND VGND VPWR VPWR _00608_ sky130_fd_sc_hd__mux2_1
Xhold2128 data_array.data1\[13\]\[37\] VGND VGND VPWR VPWR net3779 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2139 tag_array.tag0\[2\]\[14\] VGND VGND VPWR VPWR net3790 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1405 data_array.data0\[10\]\[53\] VGND VGND VPWR VPWR net3056 sky130_fd_sc_hd__dlygate4sd3_1
X_07802_ net1213 _05005_ _05009_ net1165 VGND VGND VPWR VPWR _05011_ sky130_fd_sc_hd__a22o_1
Xhold1416 data_array.data1\[3\]\[34\] VGND VGND VPWR VPWR net3067 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1427 data_array.data1\[10\]\[10\] VGND VGND VPWR VPWR net3078 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1438 data_array.data0\[6\]\[20\] VGND VGND VPWR VPWR net3089 sky130_fd_sc_hd__dlygate4sd3_1
X_05994_ data_array.rdata1\[54\] net830 net839 VGND VGND VPWR VPWR _03457_ sky130_fd_sc_hd__a21o_1
XFILLER_57_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08782_ net696 net3095 _05606_ VGND VGND VPWR VPWR _00541_ sky130_fd_sc_hd__mux2_1
XFILLER_111_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1449 data_array.data0\[2\]\[36\] VGND VGND VPWR VPWR net3100 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_940 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_4__f_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_5_4__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_07733_ data_array.data1\[1\]\[26\] net1526 net1430 data_array.data1\[2\]\[26\] VGND
+ VGND VPWR VPWR _04948_ sky130_fd_sc_hd__a22o_1
XFILLER_38_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07664_ data_array.data1\[4\]\[20\] net1419 net1325 data_array.data1\[7\]\[20\] _04884_
+ VGND VGND VPWR VPWR _04885_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_49_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09403_ net1055 net2478 net585 VGND VGND VPWR VPWR _01156_ sky130_fd_sc_hd__mux2_1
X_06615_ _03930_ _03931_ VGND VGND VPWR VPWR _00160_ sky130_fd_sc_hd__or2_1
XFILLER_164_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07595_ data_array.data1\[9\]\[14\] net1568 net1472 data_array.data1\[10\]\[14\]
+ VGND VGND VPWR VPWR _04822_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_66_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06546_ tag_array.tag1\[0\]\[7\] net1419 net1325 tag_array.tag1\[3\]\[7\] _03868_
+ VGND VGND VPWR VPWR _03869_ sky130_fd_sc_hd__a221o_1
XFILLER_80_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09334_ net1064 net3330 net406 VGND VGND VPWR VPWR _01087_ sky130_fd_sc_hd__mux2_1
XFILLER_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09265_ net718 net2243 net571 VGND VGND VPWR VPWR _01019_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06477_ tag_array.tag1\[9\]\[1\] net1542 net1446 tag_array.tag1\[10\]\[1\] VGND VGND
+ VPWR VPWR _03806_ sky130_fd_sc_hd__a22o_1
XFILLER_166_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08216_ fsm.tag_out1\[7\] net817 net809 fsm.tag_out0\[7\] _05378_ VGND VGND VPWR
+ VPWR _05379_ sky130_fd_sc_hd__a221o_2
X_09196_ net696 net3097 net629 VGND VGND VPWR VPWR _00950_ sky130_fd_sc_hd__mux2_1
XFILLER_4_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08147_ tag_array.dirty1\[1\] net1542 net1446 tag_array.dirty1\[2\] VGND VGND VPWR
+ VPWR _05324_ sky130_fd_sc_hd__a22o_1
XFILLER_101_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08078_ _05260_ _05261_ VGND VGND VPWR VPWR _00116_ sky130_fd_sc_hd__or2_1
Xclkload170 clknet_leaf_195_clk VGND VGND VPWR VPWR clkload170/X sky130_fd_sc_hd__clkbuf_8
XFILLER_105_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload181 clknet_leaf_181_clk VGND VGND VPWR VPWR clkload181/Y sky130_fd_sc_hd__clkinv_4
XFILLER_20_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload192 clknet_leaf_101_clk VGND VGND VPWR VPWR clkload192/Y sky130_fd_sc_hd__inv_8
XFILLER_134_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07029_ data_array.data0\[1\]\[26\] net1529 net1433 data_array.data0\[2\]\[26\] VGND
+ VGND VPWR VPWR _04308_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_8_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10040_ net924 net3165 net554 VGND VGND VPWR VPWR _01789_ sky130_fd_sc_hd__mux2_1
XFILLER_102_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2640 data_array.data1\[6\]\[42\] VGND VGND VPWR VPWR net4291 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_145_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2651 data_array.data0\[10\]\[44\] VGND VGND VPWR VPWR net4302 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2662 tag_array.tag0\[15\]\[18\] VGND VGND VPWR VPWR net4313 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 reset VGND VGND VPWR VPWR net1694 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold54 tag_array.valid0\[13\] VGND VGND VPWR VPWR net1705 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2673 data_array.data0\[7\]\[16\] VGND VGND VPWR VPWR net4324 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_21_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold65 tag_array.valid0\[4\] VGND VGND VPWR VPWR net1716 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_162_3470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold76 tag_array.valid1\[2\] VGND VGND VPWR VPWR net1727 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2684 tag_array.tag0\[0\]\[11\] VGND VGND VPWR VPWR net4335 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_162_3481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2695 data_array.data0\[11\]\[60\] VGND VGND VPWR VPWR net4346 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 data_array.data0\[2\]\[13\] VGND VGND VPWR VPWR net1738 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1950 data_array.data0\[10\]\[22\] VGND VGND VPWR VPWR net3601 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1961 data_array.data1\[13\]\[42\] VGND VGND VPWR VPWR net3612 sky130_fd_sc_hd__dlygate4sd3_1
X_11991_ clknet_leaf_264_clk _00799_ VGND VGND VPWR VPWR data_array.data0\[6\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1972 tag_array.tag0\[14\]\[18\] VGND VGND VPWR VPWR net3623 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 data_array.data0\[4\]\[49\] VGND VGND VPWR VPWR net1749 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1983 tag_array.tag1\[3\]\[16\] VGND VGND VPWR VPWR net3634 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13730_ clknet_leaf_255_clk _02359_ VGND VGND VPWR VPWR data_array.data1\[1\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1994 tag_array.tag1\[11\]\[3\] VGND VGND VPWR VPWR net3645 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_123_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10942_ net974 net2431 net527 VGND VGND VPWR VPWR _02687_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_123_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13661_ clknet_leaf_229_clk _02290_ VGND VGND VPWR VPWR data_array.data1\[15\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_10873_ net994 net3582 net519 VGND VGND VPWR VPWR _02618_ sky130_fd_sc_hd__mux2_1
X_12612_ clknet_leaf_106_clk _01306_ VGND VGND VPWR VPWR tag_array.tag0\[0\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_13592_ clknet_leaf_246_clk _02221_ VGND VGND VPWR VPWR data_array.data0\[9\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12543_ clknet_leaf_106_clk _01237_ VGND VGND VPWR VPWR tag_array.tag0\[11\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_129_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12474_ clknet_leaf_246_clk _01168_ VGND VGND VPWR VPWR data_array.data1\[9\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_14213_ clknet_leaf_206_clk _02842_ VGND VGND VPWR VPWR data_array.data0\[2\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11425_ clknet_leaf_50_clk _00235_ VGND VGND VPWR VPWR data_array.data0\[0\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_169_3602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_169_3613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_7 _00156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14144_ clknet_leaf_12_clk _02773_ VGND VGND VPWR VPWR data_array.data0\[1\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
X_11356_ net870 net3000 net804 VGND VGND VPWR VPWR _03099_ sky130_fd_sc_hd__mux2_1
XFILLER_126_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10307_ net2380 net935 net641 VGND VGND VPWR VPWR _02054_ sky130_fd_sc_hd__mux2_1
X_14075_ clknet_leaf_4_clk _02704_ VGND VGND VPWR VPWR data_array.data1\[6\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
X_11287_ net882 net4592 net676 VGND VGND VPWR VPWR _03030_ sky130_fd_sc_hd__mux2_1
X_13026_ clknet_leaf_260_clk _01720_ VGND VGND VPWR VPWR data_array.data0\[3\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
X_10238_ net793 net2430 net596 VGND VGND VPWR VPWR _01985_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_182_3857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1030 _05460_ VGND VGND VPWR VPWR net1030 sky130_fd_sc_hd__clkbuf_2
XFILLER_117_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1041 _05454_ VGND VGND VPWR VPWR net1041 sky130_fd_sc_hd__buf_1
X_10169_ net869 net4346 net369 VGND VGND VPWR VPWR _01917_ sky130_fd_sc_hd__mux2_1
Xfanout1052 _05448_ VGND VGND VPWR VPWR net1052 sky130_fd_sc_hd__clkbuf_2
Xfanout1063 _05444_ VGND VGND VPWR VPWR net1063 sky130_fd_sc_hd__buf_1
Xfanout1074 _05438_ VGND VGND VPWR VPWR net1074 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1085 _05432_ VGND VGND VPWR VPWR net1085 sky130_fd_sc_hd__clkbuf_2
XFILLER_82_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1096 _05426_ VGND VGND VPWR VPWR net1096 sky130_fd_sc_hd__clkbuf_2
XFILLER_47_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13928_ clknet_leaf_265_clk _02557_ VGND VGND VPWR VPWR data_array.data1\[4\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_179_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13859_ clknet_leaf_248_clk _02488_ VGND VGND VPWR VPWR data_array.data1\[3\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06400_ tag_array.tag0\[9\]\[19\] net1596 net1500 tag_array.tag0\[10\]\[19\] VGND
+ VGND VPWR VPWR _03736_ sky130_fd_sc_hd__a22o_1
X_07380_ data_array.data0\[12\]\[58\] net1357 net1263 data_array.data0\[15\]\[58\]
+ _04626_ VGND VGND VPWR VPWR _04627_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_44_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06331_ tag_array.tag0\[8\]\[13\] net1410 net1316 tag_array.tag0\[11\]\[13\] _03672_
+ VGND VGND VPWR VPWR _03673_ sky130_fd_sc_hd__a221o_1
XFILLER_176_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09050_ net1084 net2449 net410 VGND VGND VPWR VPWR _00804_ sky130_fd_sc_hd__mux2_1
X_06262_ net1172 _03605_ _03609_ net1221 VGND VGND VPWR VPWR _03611_ sky130_fd_sc_hd__a22o_1
X_08001_ _05190_ _05191_ VGND VGND VPWR VPWR _00109_ sky130_fd_sc_hd__or2_1
X_06193_ tag_array.tag0\[1\]\[0\] net1595 net1499 tag_array.tag0\[2\]\[0\] VGND VGND
+ VPWR VPWR _03548_ sky130_fd_sc_hd__a22o_1
Xhold502 data_array.data1\[2\]\[49\] VGND VGND VPWR VPWR net2153 sky130_fd_sc_hd__dlygate4sd3_1
Xhold513 data_array.data1\[0\]\[39\] VGND VGND VPWR VPWR net2164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold524 data_array.data1\[8\]\[54\] VGND VGND VPWR VPWR net2175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold535 tag_array.tag1\[10\]\[16\] VGND VGND VPWR VPWR net2186 sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 data_array.data0\[12\]\[7\] VGND VGND VPWR VPWR net2197 sky130_fd_sc_hd__dlygate4sd3_1
Xhold557 data_array.data0\[15\]\[9\] VGND VGND VPWR VPWR net2208 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold568 data_array.data0\[1\]\[48\] VGND VGND VPWR VPWR net2219 sky130_fd_sc_hd__dlygate4sd3_1
X_09952_ net1020 net3959 net371 VGND VGND VPWR VPWR _01701_ sky130_fd_sc_hd__mux2_1
XFILLER_116_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold579 data_array.data0\[2\]\[19\] VGND VGND VPWR VPWR net2230 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1010 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08903_ net895 net3821 net436 VGND VGND VPWR VPWR _00660_ sky130_fd_sc_hd__mux2_1
X_09883_ net939 net4119 net382 VGND VGND VPWR VPWR _01633_ sky130_fd_sc_hd__mux2_1
XFILLER_44_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1202 tag_array.tag1\[3\]\[0\] VGND VGND VPWR VPWR net2853 sky130_fd_sc_hd__dlygate4sd3_1
X_08834_ net1842 net909 net449 VGND VGND VPWR VPWR _00592_ sky130_fd_sc_hd__mux2_1
XFILLER_85_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1213 data_array.data1\[14\]\[0\] VGND VGND VPWR VPWR net2864 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_1079 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1224 tag_array.tag0\[7\]\[0\] VGND VGND VPWR VPWR net2875 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_170_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1235 data_array.data1\[13\]\[15\] VGND VGND VPWR VPWR net2886 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1246 tag_array.tag1\[14\]\[22\] VGND VGND VPWR VPWR net2897 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1257 data_array.data1\[6\]\[26\] VGND VGND VPWR VPWR net2908 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08765_ net762 net3630 net452 VGND VGND VPWR VPWR _00524_ sky130_fd_sc_hd__mux2_1
X_05977_ net141 net1157 _03444_ _03445_ VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__a22o_1
Xhold1268 tag_array.tag1\[7\]\[13\] VGND VGND VPWR VPWR net2919 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1279 data_array.data0\[7\]\[58\] VGND VGND VPWR VPWR net2930 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07716_ data_array.data1\[13\]\[25\] net1520 net1424 data_array.data1\[14\]\[25\]
+ VGND VGND VPWR VPWR _04932_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_140_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08696_ net1921 net740 net488 VGND VGND VPWR VPWR _00455_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_140_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07647_ net1618 _04863_ _04867_ net1192 VGND VGND VPWR VPWR _04870_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_101_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07578_ data_array.data1\[12\]\[12\] net1395 net1301 data_array.data1\[15\]\[12\]
+ _04806_ VGND VGND VPWR VPWR _04807_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_24_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_801 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09317_ net710 net4170 net544 VGND VGND VPWR VPWR _01071_ sky130_fd_sc_hd__mux2_1
X_06529_ tag_array.tag1\[12\]\[6\] net1362 net1268 tag_array.tag1\[15\]\[6\] _03852_
+ VGND VGND VPWR VPWR _03853_ sky130_fd_sc_hd__a221o_1
XFILLER_21_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09248_ net786 net4106 net568 VGND VGND VPWR VPWR _01002_ sky130_fd_sc_hd__mux2_1
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_10_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_10_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_119_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09179_ net762 net4243 net629 VGND VGND VPWR VPWR _00933_ sky130_fd_sc_hd__mux2_1
X_11210_ net935 net3910 net657 VGND VGND VPWR VPWR _02953_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12190_ clknet_leaf_181_clk _00998_ VGND VGND VPWR VPWR tag_array.tag0\[14\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_162_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11141_ net953 net3495 net543 VGND VGND VPWR VPWR _02884_ sky130_fd_sc_hd__mux2_1
XFILLER_123_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_164_3510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11072_ net2527 net972 net328 VGND VGND VPWR VPWR _02815_ sky130_fd_sc_hd__mux2_1
Xinput100 mem_rdata[10] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_1
Xinput111 mem_rdata[20] VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput122 mem_rdata[30] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_1
X_10023_ net994 net3115 net561 VGND VGND VPWR VPWR _01772_ sky130_fd_sc_hd__mux2_1
Xinput133 mem_rdata[40] VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_1
Xinput144 mem_rdata[50] VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_1
Xinput155 mem_rdata[60] VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_160_3429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2470 data_array.data0\[12\]\[39\] VGND VGND VPWR VPWR net4121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2481 data_array.data1\[3\]\[37\] VGND VGND VPWR VPWR net4132 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2492 data_array.data1\[3\]\[7\] VGND VGND VPWR VPWR net4143 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1780 data_array.data0\[10\]\[31\] VGND VGND VPWR VPWR net3431 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1791 tag_array.tag0\[15\]\[22\] VGND VGND VPWR VPWR net3442 sky130_fd_sc_hd__dlygate4sd3_1
X_11974_ clknet_leaf_39_clk _00782_ VGND VGND VPWR VPWR data_array.data0\[4\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13713_ clknet_leaf_61_clk _02342_ VGND VGND VPWR VPWR data_array.data1\[1\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_10925_ net1040 net2721 net526 VGND VGND VPWR VPWR _02670_ sky130_fd_sc_hd__mux2_1
XFILLER_147_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13644_ clknet_leaf_68_clk _02273_ VGND VGND VPWR VPWR data_array.data1\[15\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_147_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10856_ net1062 net4609 net520 VGND VGND VPWR VPWR _02601_ sky130_fd_sc_hd__mux2_1
XFILLER_60_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_862 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13575_ clknet_leaf_227_clk _02204_ VGND VGND VPWR VPWR data_array.data0\[9\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_10787_ net1979 net1082 net508 VGND VGND VPWR VPWR _02532_ sky130_fd_sc_hd__mux2_1
XFILLER_158_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12526_ clknet_leaf_137_clk _01220_ VGND VGND VPWR VPWR tag_array.tag1\[11\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12457_ clknet_leaf_58_clk _01151_ VGND VGND VPWR VPWR data_array.data1\[9\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_11408_ clknet_leaf_194_clk _00218_ VGND VGND VPWR VPWR tag_array.tag1\[7\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_10_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12388_ clknet_leaf_1_clk _01082_ VGND VGND VPWR VPWR data_array.data0\[14\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_125_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_184_3908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_184_3919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14127_ clknet_leaf_235_clk _02756_ VGND VGND VPWR VPWR data_array.data0\[1\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_154_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11339_ net938 net3832 net800 VGND VGND VPWR VPWR _03082_ sky130_fd_sc_hd__mux2_1
X_14058_ clknet_leaf_10_clk _02687_ VGND VGND VPWR VPWR data_array.data1\[6\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_86_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05900_ data_array.rdata0\[23\] net848 net1145 VGND VGND VPWR VPWR _03394_ sky130_fd_sc_hd__o21a_1
X_13009_ clknet_leaf_96_clk _01703_ VGND VGND VPWR VPWR data_array.data0\[3\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_06880_ data_array.data0\[13\]\[13\] net1553 net1457 data_array.data0\[14\]\[13\]
+ VGND VGND VPWR VPWR _04172_ sky130_fd_sc_hd__a22o_1
XFILLER_67_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_19_Left_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05831_ data_array.rdata1\[0\] net826 VGND VGND VPWR VPWR _03348_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_85_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08550_ net757 net3716 net588 VGND VGND VPWR VPWR _00318_ sky130_fd_sc_hd__mux2_1
X_05762_ fsm.tag_out1\[0\] net30 VGND VGND VPWR VPWR _03279_ sky130_fd_sc_hd__and2b_1
X_07501_ data_array.data1\[12\]\[5\] net1360 net1266 data_array.data1\[15\]\[5\] _04736_
+ VGND VGND VPWR VPWR _04737_ sky130_fd_sc_hd__a221o_1
X_08481_ net1724 net638 VGND VGND VPWR VPWR _00289_ sky130_fd_sc_hd__or2_1
X_05693_ net21 fsm.tag_out0\[21\] VGND VGND VPWR VPWR _03210_ sky130_fd_sc_hd__and2b_1
XFILLER_35_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07432_ data_array.data0\[5\]\[63\] net1556 net1460 data_array.data0\[6\]\[63\] VGND
+ VGND VPWR VPWR _04674_ sky130_fd_sc_hd__a22o_1
XFILLER_161_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07363_ _04610_ _04611_ VGND VGND VPWR VPWR _00051_ sky130_fd_sc_hd__or2_1
XFILLER_148_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Left_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09102_ net876 net3696 net413 VGND VGND VPWR VPWR _00856_ sky130_fd_sc_hd__mux2_1
X_06314_ tag_array.tag0\[5\]\[11\] net1592 net1496 tag_array.tag0\[6\]\[11\] VGND
+ VGND VPWR VPWR _03658_ sky130_fd_sc_hd__a22o_1
X_07294_ data_array.data0\[0\]\[50\] net1346 net1252 data_array.data0\[3\]\[50\] _04548_
+ VGND VGND VPWR VPWR _04549_ sky130_fd_sc_hd__a221o_1
X_09033_ net2557 net894 net420 VGND VGND VPWR VPWR _00788_ sky130_fd_sc_hd__mux2_1
X_06245_ tag_array.tag0\[4\]\[5\] net1418 net1324 tag_array.tag0\[7\]\[5\] _03594_
+ VGND VGND VPWR VPWR _03595_ sky130_fd_sc_hd__a221o_1
XFILLER_117_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold310 data_array.data1\[8\]\[35\] VGND VGND VPWR VPWR net1961 sky130_fd_sc_hd__dlygate4sd3_1
X_06176_ tag_array.valid1\[13\] net1559 net1463 tag_array.valid1\[14\] VGND VGND VPWR
+ VPWR _03532_ sky130_fd_sc_hd__a22o_1
Xhold321 data_array.data1\[0\]\[43\] VGND VGND VPWR VPWR net1972 sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 data_array.data1\[0\]\[58\] VGND VGND VPWR VPWR net1983 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold343 data_array.data1\[8\]\[55\] VGND VGND VPWR VPWR net1994 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_11_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold354 tag_array.tag1\[8\]\[10\] VGND VGND VPWR VPWR net2005 sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 data_array.data0\[4\]\[32\] VGND VGND VPWR VPWR net2016 sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 data_array.data1\[1\]\[51\] VGND VGND VPWR VPWR net2027 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold387 data_array.data1\[0\]\[62\] VGND VGND VPWR VPWR net2038 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold398 data_array.data0\[8\]\[25\] VGND VGND VPWR VPWR net2049 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout801 net803 VGND VGND VPWR VPWR net801 sky130_fd_sc_hd__clkbuf_8
X_09935_ net1088 net3224 net372 VGND VGND VPWR VPWR _01684_ sky130_fd_sc_hd__mux2_1
Xfanout812 net815 VGND VGND VPWR VPWR net812 sky130_fd_sc_hd__clkbuf_2
Xfanout823 net825 VGND VGND VPWR VPWR net823 sky130_fd_sc_hd__buf_1
Xfanout834 net835 VGND VGND VPWR VPWR net834 sky130_fd_sc_hd__buf_12
XFILLER_58_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_37_Left_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout856 net857 VGND VGND VPWR VPWR net856 sky130_fd_sc_hd__clkbuf_2
Xfanout867 _05542_ VGND VGND VPWR VPWR net867 sky130_fd_sc_hd__buf_1
X_09866_ net1006 net3200 net378 VGND VGND VPWR VPWR _01616_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_142_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1010 data_array.data1\[8\]\[19\] VGND VGND VPWR VPWR net2661 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout878 net879 VGND VGND VPWR VPWR net878 sky130_fd_sc_hd__clkbuf_2
XFILLER_133_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1021 tag_array.tag1\[9\]\[18\] VGND VGND VPWR VPWR net2672 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout889 _05530_ VGND VGND VPWR VPWR net889 sky130_fd_sc_hd__buf_1
Xhold1032 tag_array.tag0\[4\]\[15\] VGND VGND VPWR VPWR net2683 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_133_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08817_ net2964 net977 net447 VGND VGND VPWR VPWR _00575_ sky130_fd_sc_hd__mux2_1
Xhold1043 data_array.data0\[8\]\[2\] VGND VGND VPWR VPWR net2694 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1054 data_array.data1\[1\]\[25\] VGND VGND VPWR VPWR net2705 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09797_ net1022 net2946 net387 VGND VGND VPWR VPWR _01548_ sky130_fd_sc_hd__mux2_1
Xhold1065 data_array.data1\[0\]\[25\] VGND VGND VPWR VPWR net2716 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1076 tag_array.tag0\[15\]\[7\] VGND VGND VPWR VPWR net2727 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1087 data_array.data0\[6\]\[53\] VGND VGND VPWR VPWR net2738 sky130_fd_sc_hd__dlygate4sd3_1
X_08748_ net730 net2383 net465 VGND VGND VPWR VPWR _00507_ sky130_fd_sc_hd__mux2_1
XFILLER_73_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1098 tag_array.tag1\[8\]\[14\] VGND VGND VPWR VPWR net2749 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_55 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08679_ net706 net2162 net501 VGND VGND VPWR VPWR _00438_ sky130_fd_sc_hd__mux2_1
XFILLER_14_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10710_ net1887 net878 net481 VGND VGND VPWR VPWR _02455_ sky130_fd_sc_hd__mux2_1
XFILLER_159_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11690_ clknet_leaf_188_clk _00498_ VGND VGND VPWR VPWR tag_array.tag1\[15\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_46_Left_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10641_ net1802 net898 net467 VGND VGND VPWR VPWR _02386_ sky130_fd_sc_hd__mux2_1
XFILLER_139_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_3380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13360_ clknet_leaf_142_clk _01990_ VGND VGND VPWR VPWR tag_array.tag0\[2\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_10572_ net919 net4135 net461 VGND VGND VPWR VPWR _02317_ sky130_fd_sc_hd__mux2_1
XFILLER_166_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_165_Right_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12311_ clknet_leaf_187_clk _01069_ VGND VGND VPWR VPWR tag_array.tag1\[12\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_153_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13291_ clknet_leaf_227_clk _01921_ VGND VGND VPWR VPWR data_array.data0\[10\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12242_ clknet_leaf_184_clk _00172_ VGND VGND VPWR VPWR fsm.tag_out1\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12173_ clknet_leaf_144_clk _00981_ VGND VGND VPWR VPWR tag_array.tag0\[14\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_131_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_55_Left_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11124_ net1021 net4003 net543 VGND VGND VPWR VPWR _02867_ sky130_fd_sc_hd__mux2_1
XFILLER_96_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_992 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11055_ net2632 net1042 net331 VGND VGND VPWR VPWR _02798_ sky130_fd_sc_hd__mux2_1
XFILLER_122_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10006_ net1063 net3085 net562 VGND VGND VPWR VPWR _01755_ sky130_fd_sc_hd__mux2_1
XFILLER_37_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11957_ clknet_leaf_34_clk _00765_ VGND VGND VPWR VPWR data_array.data0\[4\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_91_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_177_3756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_177_3767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10908_ net1110 net3609 net529 VGND VGND VPWR VPWR _02653_ sky130_fd_sc_hd__mux2_1
X_11888_ clknet_leaf_247_clk _00696_ VGND VGND VPWR VPWR data_array.data0\[5\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13627_ clknet_leaf_223_clk _02256_ VGND VGND VPWR VPWR data_array.data0\[9\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10839_ net1981 net875 net507 VGND VGND VPWR VPWR _02584_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_1053 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13558_ clknet_leaf_17_clk _02187_ VGND VGND VPWR VPWR data_array.data1\[0\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_132_Right_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12509_ clknet_leaf_210_clk _01203_ VGND VGND VPWR VPWR data_array.data1\[9\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
X_13489_ clknet_leaf_171_clk _02119_ VGND VGND VPWR VPWR tag_array.tag0\[15\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_66_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06030_ _03476_ net1131 VGND VGND VPWR VPWR _03480_ sky130_fd_sc_hd__or2_4
XFILLER_145_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07981_ data_array.data1\[12\]\[49\] net1381 net1287 data_array.data1\[15\]\[49\]
+ _05172_ VGND VGND VPWR VPWR _05173_ sky130_fd_sc_hd__a221o_1
XFILLER_86_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09720_ net709 net2600 net611 VGND VGND VPWR VPWR _01472_ sky130_fd_sc_hd__mux2_1
X_06932_ net1190 _04213_ _04217_ net1616 VGND VGND VPWR VPWR _04220_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09651_ net784 net4265 net612 VGND VGND VPWR VPWR _01403_ sky130_fd_sc_hd__mux2_1
X_06863_ data_array.data0\[12\]\[11\] net1383 net1289 data_array.data0\[15\]\[11\]
+ _04156_ VGND VGND VPWR VPWR _04157_ sky130_fd_sc_hd__a221o_1
X_08602_ net714 net4383 net534 VGND VGND VPWR VPWR _00361_ sky130_fd_sc_hd__mux2_1
X_05814_ _03173_ _03187_ _03188_ _03218_ VGND VGND VPWR VPWR _03331_ sky130_fd_sc_hd__or4_1
X_09582_ net1022 net4466 net395 VGND VGND VPWR VPWR _01334_ sky130_fd_sc_hd__mux2_1
X_06794_ data_array.data0\[1\]\[5\] net1546 net1450 data_array.data0\[2\]\[5\] VGND
+ VGND VPWR VPWR _04094_ sky130_fd_sc_hd__a22o_1
X_08533_ _05558_ net815 VGND VGND VPWR VPWR _05593_ sky130_fd_sc_hd__nand2b_4
XFILLER_36_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05745_ _03258_ _03259_ _03260_ _03261_ VGND VGND VPWR VPWR _03262_ sky130_fd_sc_hd__or4_1
X_08464_ net1126 _05545_ VGND VGND VPWR VPWR _05546_ sky130_fd_sc_hd__and2_1
X_05676_ fsm.tag_out0\[20\] net20 VGND VGND VPWR VPWR _03193_ sky130_fd_sc_hd__and2b_1
X_07415_ data_array.data0\[4\]\[61\] net1357 net1263 data_array.data0\[7\]\[61\] _04658_
+ VGND VGND VPWR VPWR _04659_ sky130_fd_sc_hd__a221o_1
X_08395_ net1129 _05499_ VGND VGND VPWR VPWR _05500_ sky130_fd_sc_hd__and2_1
XFILLER_177_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07346_ data_array.data0\[9\]\[55\] net1534 net1438 data_array.data0\[10\]\[55\]
+ VGND VGND VPWR VPWR _04596_ sky130_fd_sc_hd__a22o_1
XFILLER_148_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07277_ data_array.data0\[12\]\[49\] net1380 net1286 data_array.data0\[15\]\[49\]
+ _04532_ VGND VGND VPWR VPWR _04533_ sky130_fd_sc_hd__a221o_1
XFILLER_128_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09016_ net2078 net962 net420 VGND VGND VPWR VPWR _00771_ sky130_fd_sc_hd__mux2_1
X_06228_ net1200 _03573_ _03577_ net1626 VGND VGND VPWR VPWR _03580_ sky130_fd_sc_hd__a22o_1
XFILLER_136_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06159_ net26 net27 VGND VGND VPWR VPWR _03516_ sky130_fd_sc_hd__nand2_1
Xhold140 data_array.data0\[2\]\[9\] VGND VGND VPWR VPWR net1791 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 data_array.data1\[1\]\[53\] VGND VGND VPWR VPWR net1802 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold162 data_array.data1\[2\]\[61\] VGND VGND VPWR VPWR net1813 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 tag_array.tag1\[2\]\[5\] VGND VGND VPWR VPWR net1824 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_160_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold184 data_array.data1\[8\]\[50\] VGND VGND VPWR VPWR net1835 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 tag_array.tag1\[8\]\[0\] VGND VGND VPWR VPWR net1846 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout1607 net1609 VGND VGND VPWR VPWR net1607 sky130_fd_sc_hd__clkbuf_4
Xfanout620 _05569_ VGND VGND VPWR VPWR net620 sky130_fd_sc_hd__buf_4
Xfanout1618 net1620 VGND VGND VPWR VPWR net1618 sky130_fd_sc_hd__buf_4
Xfanout1629 _03506_ VGND VGND VPWR VPWR net1629 sky130_fd_sc_hd__buf_4
Xfanout631 net632 VGND VGND VPWR VPWR net631 sky130_fd_sc_hd__buf_4
XFILLER_120_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout642 net643 VGND VGND VPWR VPWR net642 sky130_fd_sc_hd__buf_4
X_09918_ net736 net2437 net602 VGND VGND VPWR VPWR _01668_ sky130_fd_sc_hd__mux2_1
Xfanout653 net654 VGND VGND VPWR VPWR net653 sky130_fd_sc_hd__buf_2
Xfanout664 net665 VGND VGND VPWR VPWR net664 sky130_fd_sc_hd__buf_4
Xfanout675 net676 VGND VGND VPWR VPWR net675 sky130_fd_sc_hd__clkbuf_8
XFILLER_19_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout686 net690 VGND VGND VPWR VPWR net686 sky130_fd_sc_hd__buf_4
X_09849_ net1072 net2675 net383 VGND VGND VPWR VPWR _01599_ sky130_fd_sc_hd__mux2_1
XFILLER_74_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout697 _05413_ VGND VGND VPWR VPWR net697 sky130_fd_sc_hd__clkbuf_2
XFILLER_92_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12860_ clknet_leaf_33_clk _01554_ VGND VGND VPWR VPWR data_array.data0\[12\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_170_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11811_ clknet_leaf_206_clk _00619_ VGND VGND VPWR VPWR data_array.data0\[7\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_159_3420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ clknet_leaf_141_clk _01485_ VGND VGND VPWR VPWR tag_array.tag1\[10\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11742_ clknet_leaf_16_clk _00550_ VGND VGND VPWR VPWR data_array.data0\[8\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_155_3339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461_ clknet_leaf_26_clk _03084_ VGND VGND VPWR VPWR data_array.data1\[7\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11673_ clknet_leaf_168_clk _00481_ VGND VGND VPWR VPWR tag_array.tag1\[1\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_13412_ clknet_leaf_258_clk _02042_ VGND VGND VPWR VPWR data_array.data1\[8\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_12_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10624_ net1942 net965 net472 VGND VGND VPWR VPWR _02369_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14392_ clknet_leaf_88_clk _03015_ VGND VGND VPWR VPWR data_array.data1\[10\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_172_3675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13343_ clknet_leaf_223_clk _01973_ VGND VGND VPWR VPWR data_array.data0\[10\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
X_10555_ net985 net2507 net460 VGND VGND VPWR VPWR _02300_ sky130_fd_sc_hd__mux2_1
XFILLER_139_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_133_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13274_ clknet_leaf_91_clk _01904_ VGND VGND VPWR VPWR data_array.data0\[11\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
X_10486_ net1002 net4287 net347 VGND VGND VPWR VPWR _02231_ sky130_fd_sc_hd__mux2_1
XFILLER_52_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12225_ clknet_leaf_145_clk _00178_ VGND VGND VPWR VPWR fsm.tag_out1\[7\] sky130_fd_sc_hd__dfxtp_1
X_12156_ clknet_leaf_145_clk _00964_ VGND VGND VPWR VPWR tag_array.tag0\[13\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_151_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11107_ net1091 net3090 net545 VGND VGND VPWR VPWR _02850_ sky130_fd_sc_hd__mux2_1
XFILLER_1_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12087_ clknet_leaf_75_clk _00895_ VGND VGND VPWR VPWR data_array.data1\[14\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_34_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11038_ net2199 net1108 net332 VGND VGND VPWR VPWR _02781_ sky130_fd_sc_hd__mux2_1
XFILLER_76_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_179_3807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_334 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_1071 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12989_ clknet_leaf_72_clk _01683_ VGND VGND VPWR VPWR data_array.data0\[3\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_178_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_940 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_180_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_180_clk
+ sky130_fd_sc_hd__clkbuf_8
X_07200_ data_array.data0\[8\]\[42\] net1386 net1292 data_array.data0\[11\]\[42\]
+ _04462_ VGND VGND VPWR VPWR _04463_ sky130_fd_sc_hd__a221o_1
XFILLER_32_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08180_ net1644 net33 net4624 VGND VGND VPWR VPWR _00184_ sky130_fd_sc_hd__o21a_1
XFILLER_118_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07131_ net1166 _04395_ _04399_ net1214 VGND VGND VPWR VPWR _04401_ sky130_fd_sc_hd__a22o_1
XFILLER_146_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07062_ data_array.data0\[5\]\[29\] net1570 net1474 data_array.data0\[6\]\[29\] VGND
+ VGND VPWR VPWR _04338_ sky130_fd_sc_hd__a22o_1
Xoutput201 net201 VGND VGND VPWR VPWR cpu_rdata[42] sky130_fd_sc_hd__buf_6
XFILLER_161_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06013_ net155 net1157 _03468_ _03469_ VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__a22o_1
Xoutput212 net212 VGND VGND VPWR VPWR cpu_rdata[52] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_93_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput223 net223 VGND VGND VPWR VPWR cpu_rdata[62] sky130_fd_sc_hd__buf_2
XFILLER_161_659 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput234 net234 VGND VGND VPWR VPWR mem_addr[13] sky130_fd_sc_hd__buf_2
Xoutput245 net245 VGND VGND VPWR VPWR mem_addr[23] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput256 net256 VGND VGND VPWR VPWR mem_addr[4] sky130_fd_sc_hd__buf_2
Xoutput267 net267 VGND VGND VPWR VPWR mem_wdata[13] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput278 net278 VGND VGND VPWR VPWR mem_wdata[23] sky130_fd_sc_hd__buf_2
Xoutput289 net289 VGND VGND VPWR VPWR mem_wdata[33] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_71_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07964_ data_array.data1\[1\]\[47\] net1588 net1492 data_array.data1\[2\]\[47\] VGND
+ VGND VPWR VPWR _05158_ sky130_fd_sc_hd__a22o_1
XFILLER_68_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09703_ net776 net4369 net609 VGND VGND VPWR VPWR _01455_ sky130_fd_sc_hd__mux2_1
X_06915_ data_array.data0\[5\]\[16\] net1547 net1451 data_array.data0\[6\]\[16\] VGND
+ VGND VPWR VPWR _04204_ sky130_fd_sc_hd__a22o_1
XFILLER_114_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07895_ data_array.data1\[4\]\[41\] net1335 net1241 data_array.data1\[7\]\[41\] _05094_
+ VGND VGND VPWR VPWR _05095_ sky130_fd_sc_hd__a221o_1
X_09634_ net752 net3485 net616 VGND VGND VPWR VPWR _01386_ sky130_fd_sc_hd__mux2_1
XFILLER_67_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06846_ _04140_ _04141_ VGND VGND VPWR VPWR _00063_ sky130_fd_sc_hd__or2_1
XFILLER_167_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09565_ net1089 net3042 net396 VGND VGND VPWR VPWR _01317_ sky130_fd_sc_hd__mux2_1
X_06777_ data_array.data0\[0\]\[3\] net1377 net1283 data_array.data0\[3\]\[3\] _04078_
+ VGND VGND VPWR VPWR _04079_ sky130_fd_sc_hd__a221o_1
XFILLER_71_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08516_ net822 net811 net854 _05580_ VGND VGND VPWR VPWR _05582_ sky130_fd_sc_hd__or4b_1
XFILLER_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05728_ net19 fsm.tag_out1\[19\] VGND VGND VPWR VPWR _03245_ sky130_fd_sc_hd__xor2_1
X_09496_ net744 net2733 net624 VGND VGND VPWR VPWR _01249_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_137_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_776 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08447_ net2278 net880 net690 VGND VGND VPWR VPWR _00278_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_171_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_171_clk
+ sky130_fd_sc_hd__clkbuf_8
X_05659_ _03172_ _03173_ _03174_ _03175_ VGND VGND VPWR VPWR _03176_ sky130_fd_sc_hd__or4_1
XFILLER_184_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08378_ net3082 net972 net686 VGND VGND VPWR VPWR _00255_ sky130_fd_sc_hd__mux2_1
X_07329_ net1215 _04575_ _04579_ net1167 VGND VGND VPWR VPWR _04581_ sky130_fd_sc_hd__a22o_1
XFILLER_109_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10340_ net739 net2752 net593 VGND VGND VPWR VPWR _02087_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10271_ net2365 net1078 net635 VGND VGND VPWR VPWR _02018_ sky130_fd_sc_hd__mux2_1
XFILLER_180_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12010_ clknet_leaf_126_clk _00818_ VGND VGND VPWR VPWR data_array.data0\[6\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1404 net1406 VGND VGND VPWR VPWR net1404 sky130_fd_sc_hd__clkbuf_4
XFILLER_105_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1415 net1416 VGND VGND VPWR VPWR net1415 sky130_fd_sc_hd__clkbuf_4
Xfanout1426 net1428 VGND VGND VPWR VPWR net1426 sky130_fd_sc_hd__clkbuf_4
Xfanout1437 net1447 VGND VGND VPWR VPWR net1437 sky130_fd_sc_hd__buf_2
Xfanout1448 net1450 VGND VGND VPWR VPWR net1448 sky130_fd_sc_hd__clkbuf_4
Xfanout450 _05606_ VGND VGND VPWR VPWR net450 sky130_fd_sc_hd__buf_4
Xfanout461 net465 VGND VGND VPWR VPWR net461 sky130_fd_sc_hd__buf_4
XFILLER_48_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1459 net1461 VGND VGND VPWR VPWR net1459 sky130_fd_sc_hd__clkbuf_4
XFILLER_150_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout472 net474 VGND VGND VPWR VPWR net472 sky130_fd_sc_hd__clkbuf_8
XFILLER_63_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13961_ clknet_leaf_266_clk _02590_ VGND VGND VPWR VPWR data_array.data1\[5\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout483 net486 VGND VGND VPWR VPWR net483 sky130_fd_sc_hd__clkbuf_8
XFILLER_58_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout494 net495 VGND VGND VPWR VPWR net494 sky130_fd_sc_hd__clkbuf_8
XFILLER_86_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12912_ clknet_leaf_222_clk _01606_ VGND VGND VPWR VPWR data_array.data0\[13\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_13892_ clknet_leaf_120_clk _02521_ VGND VGND VPWR VPWR data_array.data1\[3\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_126_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12843_ clknet_leaf_45_clk _01537_ VGND VGND VPWR VPWR data_array.data0\[12\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_17_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_174_3704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ clknet_leaf_109_clk _01468_ VGND VGND VPWR VPWR tag_array.tag0\[6\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_11725_ clknet_leaf_157_clk _00533_ VGND VGND VPWR VPWR tag_array.tag0\[9\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_162_clk clknet_5_28__leaf_clk VGND VGND VPWR VPWR clknet_leaf_162_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_159_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14444_ clknet_leaf_30_clk _03067_ VGND VGND VPWR VPWR data_array.data1\[7\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_11656_ clknet_leaf_197_clk _00464_ VGND VGND VPWR VPWR tag_array.tag1\[2\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_80_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_1053 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10607_ net1873 net1034 net472 VGND VGND VPWR VPWR _02352_ sky130_fd_sc_hd__mux2_1
X_14375_ clknet_leaf_268_clk _02998_ VGND VGND VPWR VPWR data_array.data1\[10\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_11587_ clknet_leaf_191_clk _00395_ VGND VGND VPWR VPWR tag_array.tag1\[4\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13326_ clknet_leaf_243_clk _01956_ VGND VGND VPWR VPWR data_array.data0\[10\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_171_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold909 data_array.data1\[8\]\[63\] VGND VGND VPWR VPWR net2560 sky130_fd_sc_hd__dlygate4sd3_1
X_10538_ net1055 net2544 net460 VGND VGND VPWR VPWR _02283_ sky130_fd_sc_hd__mux2_1
XFILLER_143_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13257_ clknet_leaf_71_clk _01887_ VGND VGND VPWR VPWR data_array.data0\[11\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_170_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10469_ net1069 net3694 net350 VGND VGND VPWR VPWR _02214_ sky130_fd_sc_hd__mux2_1
X_12208_ clknet_leaf_151_clk _00137_ VGND VGND VPWR VPWR fsm.tag_out0\[15\] sky130_fd_sc_hd__dfxtp_1
X_13188_ clknet_leaf_267_clk _00081_ VGND VGND VPWR VPWR data_array.rdata1\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_9_1038 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12139_ clknet_leaf_155_clk _00947_ VGND VGND VPWR VPWR tag_array.tag0\[12\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_32_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1609 tag_array.tag0\[8\]\[5\] VGND VGND VPWR VPWR net3260 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_824 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06700_ tag_array.tag1\[0\]\[21\] net1403 net1309 tag_array.tag1\[3\]\[21\] _04008_
+ VGND VGND VPWR VPWR _04009_ sky130_fd_sc_hd__a221o_1
X_07680_ net1621 _04893_ _04897_ net1198 VGND VGND VPWR VPWR _04900_ sky130_fd_sc_hd__a22o_1
XFILLER_37_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_356 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06631_ tag_array.tag1\[13\]\[15\] net1594 net1498 tag_array.tag1\[14\]\[15\] VGND
+ VGND VPWR VPWR _03946_ sky130_fd_sc_hd__a22o_1
XFILLER_80_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09350_ net1002 net4375 net405 VGND VGND VPWR VPWR _01103_ sky130_fd_sc_hd__mux2_1
X_06562_ tag_array.tag1\[8\]\[9\] net1418 net1324 tag_array.tag1\[11\]\[9\] _03882_
+ VGND VGND VPWR VPWR _03883_ sky130_fd_sc_hd__a221o_1
X_08301_ net162 net97 net1640 VGND VGND VPWR VPWR _05437_ sky130_fd_sc_hd__mux2_1
X_09281_ net756 net4006 net564 VGND VGND VPWR VPWR _01035_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06493_ net1175 _03815_ _03819_ net1223 VGND VGND VPWR VPWR _03821_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_153_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_153_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_47_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08232_ net743 net4456 net805 VGND VGND VPWR VPWR _00208_ sky130_fd_sc_hd__mux2_1
XFILLER_21_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08163_ tag_array.dirty0\[4\] net1403 net1309 tag_array.dirty0\[7\] _05338_ VGND
+ VGND VPWR VPWR _05339_ sky130_fd_sc_hd__a221o_1
XFILLER_158_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07114_ data_array.data0\[4\]\[34\] net1340 net1246 data_array.data0\[7\]\[34\] _04384_
+ VGND VGND VPWR VPWR _04385_ sky130_fd_sc_hd__a221o_1
XFILLER_119_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08094_ data_array.data1\[13\]\[59\] net1572 net1476 data_array.data1\[14\]\[59\]
+ VGND VGND VPWR VPWR _05276_ sky130_fd_sc_hd__a22o_1
XFILLER_118_166 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload60 clknet_leaf_26_clk VGND VGND VPWR VPWR clkload60/Y sky130_fd_sc_hd__inv_6
Xclkload71 clknet_leaf_237_clk VGND VGND VPWR VPWR clkload71/Y sky130_fd_sc_hd__clkinv_8
X_07045_ data_array.data0\[9\]\[28\] net1542 net1446 data_array.data0\[10\]\[28\]
+ VGND VGND VPWR VPWR _04322_ sky130_fd_sc_hd__a22o_1
Xclkload82 clknet_leaf_42_clk VGND VGND VPWR VPWR clkload82/Y sky130_fd_sc_hd__clkinv_4
XFILLER_162_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload93 clknet_leaf_66_clk VGND VGND VPWR VPWR clkload93/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2800 data_array.data1\[3\]\[14\] VGND VGND VPWR VPWR net4451 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2811 data_array.data1\[12\]\[32\] VGND VGND VPWR VPWR net4462 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_47_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08996_ net1882 net1042 net420 VGND VGND VPWR VPWR _00751_ sky130_fd_sc_hd__mux2_1
Xhold2822 data_array.data0\[5\]\[21\] VGND VGND VPWR VPWR net4473 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2833 data_array.data0\[15\]\[49\] VGND VGND VPWR VPWR net4484 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_10_Left_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2844 tag_array.tag1\[5\]\[24\] VGND VGND VPWR VPWR net4495 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2855 data_array.data0\[9\]\[55\] VGND VGND VPWR VPWR net4506 sky130_fd_sc_hd__dlygate4sd3_1
X_07947_ data_array.data1\[9\]\[46\] net1527 net1431 data_array.data1\[10\]\[46\]
+ VGND VGND VPWR VPWR _05142_ sky130_fd_sc_hd__a22o_1
XFILLER_130_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2866 tag_array.tag0\[4\]\[7\] VGND VGND VPWR VPWR net4517 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2877 data_array.data1\[6\]\[46\] VGND VGND VPWR VPWR net4528 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2888 tag_array.tag1\[9\]\[24\] VGND VGND VPWR VPWR net4539 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2899 tag_array.tag0\[1\]\[2\] VGND VGND VPWR VPWR net4550 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07878_ net1619 _05073_ _05077_ net1193 VGND VGND VPWR VPWR _05080_ sky130_fd_sc_hd__a22o_1
XFILLER_83_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09617_ net880 net4317 net397 VGND VGND VPWR VPWR _01369_ sky130_fd_sc_hd__mux2_1
XFILLER_43_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06829_ data_array.data0\[9\]\[8\] net1536 net1440 data_array.data0\[10\]\[8\] VGND
+ VGND VPWR VPWR _04126_ sky130_fd_sc_hd__a22o_1
X_09548_ net735 net2914 net618 VGND VGND VPWR VPWR _01301_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_104_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09479_ net711 net4035 net651 VGND VGND VPWR VPWR _01232_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_121_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_144_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_144_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_54_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11510_ clknet_leaf_141_clk _00318_ VGND VGND VPWR VPWR tag_array.tag1\[9\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_141_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12490_ clknet_leaf_88_clk _01184_ VGND VGND VPWR VPWR data_array.data1\[9\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11441_ clknet_leaf_71_clk _00251_ VGND VGND VPWR VPWR data_array.data0\[0\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14160_ clknet_leaf_14_clk _02789_ VGND VGND VPWR VPWR data_array.data0\[2\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_164_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11372_ net1647 net3074 net625 VGND VGND VPWR VPWR _03115_ sky130_fd_sc_hd__mux2_1
XFILLER_125_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13111_ clknet_leaf_121_clk _01805_ VGND VGND VPWR VPWR data_array.data1\[13\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_166_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10323_ net2075 net871 net642 VGND VGND VPWR VPWR _02070_ sky130_fd_sc_hd__mux2_1
XFILLER_4_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14091_ clknet_leaf_48_clk _02720_ VGND VGND VPWR VPWR data_array.data0\[1\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13042_ clknet_leaf_236_clk _01736_ VGND VGND VPWR VPWR data_array.data0\[3\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
X_10254_ net726 net3156 net597 VGND VGND VPWR VPWR _02001_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_167_3563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_3574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1201 net1212 VGND VGND VPWR VPWR net1201 sky130_fd_sc_hd__buf_2
XFILLER_182_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1212 _03522_ VGND VGND VPWR VPWR net1212 sky130_fd_sc_hd__buf_4
XFILLER_59_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1223 _03518_ VGND VGND VPWR VPWR net1223 sky130_fd_sc_hd__buf_4
X_10185_ net1065 net4081 net358 VGND VGND VPWR VPWR _01932_ sky130_fd_sc_hd__mux2_1
XFILLER_132_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1234 _03518_ VGND VGND VPWR VPWR net1234 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_128_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1245 net1282 VGND VGND VPWR VPWR net1245 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_128_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1256 net1258 VGND VGND VPWR VPWR net1256 sky130_fd_sc_hd__clkbuf_4
XFILLER_94_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1267 net1269 VGND VGND VPWR VPWR net1267 sky130_fd_sc_hd__clkbuf_4
Xfanout1278 net1281 VGND VGND VPWR VPWR net1278 sky130_fd_sc_hd__clkbuf_4
XFILLER_19_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1289 net1306 VGND VGND VPWR VPWR net1289 sky130_fd_sc_hd__clkbuf_2
X_13944_ clknet_leaf_73_clk _02573_ VGND VGND VPWR VPWR data_array.data1\[4\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13875_ clknet_leaf_36_clk _02504_ VGND VGND VPWR VPWR data_array.data1\[3\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12826_ clknet_leaf_103_clk _01520_ VGND VGND VPWR VPWR tag_array.tag1\[0\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12757_ clknet_leaf_105_clk _01451_ VGND VGND VPWR VPWR tag_array.tag0\[6\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_135_clk clknet_5_31__leaf_clk VGND VGND VPWR VPWR clknet_leaf_135_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_43_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11708_ clknet_leaf_187_clk _00516_ VGND VGND VPWR VPWR tag_array.tag1\[15\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_147_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12688_ clknet_leaf_180_clk _01382_ VGND VGND VPWR VPWR tag_array.tag0\[8\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_175_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14427_ clknet_leaf_35_clk _03050_ VGND VGND VPWR VPWR data_array.data1\[7\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_11639_ clknet_leaf_135_clk _00447_ VGND VGND VPWR VPWR tag_array.tag1\[2\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14358_ clknet_leaf_18_clk _02981_ VGND VGND VPWR VPWR data_array.data1\[10\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_156_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold706 tag_array.tag1\[0\]\[6\] VGND VGND VPWR VPWR net2357 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_157_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold717 data_array.data0\[1\]\[18\] VGND VGND VPWR VPWR net2368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold728 data_array.data1\[10\]\[46\] VGND VGND VPWR VPWR net2379 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13309_ clknet_leaf_48_clk _01939_ VGND VGND VPWR VPWR data_array.data0\[10\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_90_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold739 data_array.data1\[12\]\[37\] VGND VGND VPWR VPWR net2390 sky130_fd_sc_hd__dlygate4sd3_1
X_14289_ clknet_leaf_57_clk _02918_ VGND VGND VPWR VPWR data_array.data1\[11\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_170_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2107 tag_array.tag1\[10\]\[9\] VGND VGND VPWR VPWR net3758 sky130_fd_sc_hd__dlygate4sd3_1
X_08850_ net1106 net4615 net434 VGND VGND VPWR VPWR _00607_ sky130_fd_sc_hd__mux2_1
Xhold2118 data_array.data1\[3\]\[27\] VGND VGND VPWR VPWR net3769 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2129 data_array.data1\[12\]\[55\] VGND VGND VPWR VPWR net3780 sky130_fd_sc_hd__dlygate4sd3_1
X_07801_ net1188 _05003_ _05007_ net1614 VGND VGND VPWR VPWR _05010_ sky130_fd_sc_hd__a22o_1
Xhold1406 tag_array.tag1\[14\]\[12\] VGND VGND VPWR VPWR net3057 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1417 data_array.data1\[8\]\[20\] VGND VGND VPWR VPWR net3068 sky130_fd_sc_hd__dlygate4sd3_1
X_08781_ net698 net4250 net451 VGND VGND VPWR VPWR _00540_ sky130_fd_sc_hd__mux2_1
X_05993_ data_array.rdata0\[54\] net848 net1144 VGND VGND VPWR VPWR _03456_ sky130_fd_sc_hd__o21a_1
XFILLER_38_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1428 tag_array.tag0\[6\]\[0\] VGND VGND VPWR VPWR net3079 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1439 data_array.data1\[12\]\[5\] VGND VGND VPWR VPWR net3090 sky130_fd_sc_hd__dlygate4sd3_1
X_07732_ data_array.data1\[12\]\[26\] net1335 net1241 data_array.data1\[15\]\[26\]
+ _04946_ VGND VGND VPWR VPWR _04947_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_88_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07663_ data_array.data1\[5\]\[20\] net1610 net1514 data_array.data1\[6\]\[20\] VGND
+ VGND VPWR VPWR _04884_ sky130_fd_sc_hd__a22o_1
XFILLER_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09402_ net1057 net2434 net582 VGND VGND VPWR VPWR _01155_ sky130_fd_sc_hd__mux2_1
XFILLER_19_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06614_ net1185 _03925_ _03929_ net1233 VGND VGND VPWR VPWR _03931_ sky130_fd_sc_hd__a22o_1
XFILLER_92_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07594_ _04820_ _04821_ VGND VGND VPWR VPWR _00068_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_66_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09333_ net1068 net2258 net408 VGND VGND VPWR VPWR _01086_ sky130_fd_sc_hd__mux2_1
X_06545_ tag_array.tag1\[1\]\[7\] net1610 net1514 tag_array.tag1\[2\]\[7\] VGND VGND
+ VPWR VPWR _03868_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_126_clk clknet_5_27__leaf_clk VGND VGND VPWR VPWR clknet_leaf_126_clk
+ sky130_fd_sc_hd__clkbuf_8
X_09264_ net724 net2336 net576 VGND VGND VPWR VPWR _01018_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06476_ tag_array.tag1\[4\]\[1\] net1401 net1307 tag_array.tag1\[7\]\[1\] _03804_
+ VGND VGND VPWR VPWR _03805_ sky130_fd_sc_hd__a221o_1
XFILLER_178_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08215_ net1650 net1164 net6 VGND VGND VPWR VPWR _05378_ sky130_fd_sc_hd__and3_1
XFILLER_53_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09195_ net699 net4213 net628 VGND VGND VPWR VPWR _00949_ sky130_fd_sc_hd__mux2_1
X_08146_ tag_array.dirty1\[12\] net1384 net1290 tag_array.dirty1\[15\] _05322_ VGND
+ VGND VPWR VPWR _05323_ sky130_fd_sc_hd__a221o_1
XFILLER_107_637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08077_ net1215 _05255_ _05259_ net1166 VGND VGND VPWR VPWR _05261_ sky130_fd_sc_hd__a22o_1
Xclkload160 clknet_leaf_173_clk VGND VGND VPWR VPWR clkload160/Y sky130_fd_sc_hd__inv_6
XFILLER_134_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload171 clknet_leaf_196_clk VGND VGND VPWR VPWR clkload171/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_84_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload182 clknet_leaf_183_clk VGND VGND VPWR VPWR clkload182/Y sky130_fd_sc_hd__inv_6
XFILLER_161_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload193 clknet_leaf_102_clk VGND VGND VPWR VPWR clkload193/Y sky130_fd_sc_hd__clkinv_4
X_07028_ data_array.data0\[12\]\[26\] net1337 net1243 data_array.data0\[15\]\[26\]
+ _04306_ VGND VGND VPWR VPWR _04307_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_8_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2630 data_array.data1\[12\]\[54\] VGND VGND VPWR VPWR net4281 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2641 data_array.data1\[7\]\[1\] VGND VGND VPWR VPWR net4292 sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ net2739 net1108 net421 VGND VGND VPWR VPWR _00734_ sky130_fd_sc_hd__mux2_1
Xhold44 tag_array.valid1\[6\] VGND VGND VPWR VPWR net1695 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2652 tag_array.tag0\[3\]\[23\] VGND VGND VPWR VPWR net4303 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2663 data_array.data1\[10\]\[53\] VGND VGND VPWR VPWR net4314 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 tag_array.valid0\[10\] VGND VGND VPWR VPWR net1706 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2674 data_array.data0\[14\]\[6\] VGND VGND VPWR VPWR net4325 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_162_3471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2685 data_array.data1\[7\]\[48\] VGND VGND VPWR VPWR net4336 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1940 data_array.data0\[9\]\[50\] VGND VGND VPWR VPWR net3591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 tag_array.valid0\[3\] VGND VGND VPWR VPWR net1717 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold77 tag_array.valid1\[0\] VGND VGND VPWR VPWR net1728 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1951 tag_array.tag0\[7\]\[20\] VGND VGND VPWR VPWR net3602 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11990_ clknet_leaf_230_clk _00798_ VGND VGND VPWR VPWR data_array.data0\[6\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2696 data_array.data0\[6\]\[14\] VGND VGND VPWR VPWR net4347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 data_array.data0\[1\]\[49\] VGND VGND VPWR VPWR net1739 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_60_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1962 tag_array.tag1\[10\]\[2\] VGND VGND VPWR VPWR net3613 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 data_array.data0\[0\]\[49\] VGND VGND VPWR VPWR net1750 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1973 data_array.data1\[5\]\[56\] VGND VGND VPWR VPWR net3624 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1984 data_array.data1\[15\]\[20\] VGND VGND VPWR VPWR net3635 sky130_fd_sc_hd__dlygate4sd3_1
X_10941_ net978 net3571 net533 VGND VGND VPWR VPWR _02686_ sky130_fd_sc_hd__mux2_1
Xhold1995 data_array.data0\[9\]\[51\] VGND VGND VPWR VPWR net3646 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_123_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13660_ clknet_leaf_130_clk _02289_ VGND VGND VPWR VPWR data_array.data1\[15\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_10872_ net996 net3478 net518 VGND VGND VPWR VPWR _02617_ sky130_fd_sc_hd__mux2_1
XFILLER_44_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12611_ clknet_leaf_183_clk _01305_ VGND VGND VPWR VPWR tag_array.tag0\[0\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_117_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_117_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13591_ clknet_leaf_224_clk _02220_ VGND VGND VPWR VPWR data_array.data0\[9\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_43_189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12542_ clknet_leaf_188_clk _01236_ VGND VGND VPWR VPWR tag_array.tag1\[11\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12473_ clknet_leaf_267_clk _01167_ VGND VGND VPWR VPWR data_array.data1\[9\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14212_ clknet_leaf_114_clk _02841_ VGND VGND VPWR VPWR data_array.data0\[2\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11424_ clknet_leaf_206_clk _00234_ VGND VGND VPWR VPWR data_array.data0\[0\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_172_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_169_3603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_169_3614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_8 _00156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14143_ clknet_leaf_14_clk _02772_ VGND VGND VPWR VPWR data_array.data0\[1\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
X_11355_ net875 net4046 net800 VGND VGND VPWR VPWR _03098_ sky130_fd_sc_hd__mux2_1
XFILLER_4_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10306_ net1865 net938 net639 VGND VGND VPWR VPWR _02053_ sky130_fd_sc_hd__mux2_1
X_14074_ clknet_leaf_245_clk _02703_ VGND VGND VPWR VPWR data_array.data1\[6\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
X_11286_ net886 net2938 net675 VGND VGND VPWR VPWR _03029_ sky130_fd_sc_hd__mux2_1
XFILLER_141_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13025_ clknet_leaf_125_clk _01719_ VGND VGND VPWR VPWR data_array.data0\[3\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_112_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10237_ net857 net4541 net357 VGND VGND VPWR VPWR _01984_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_182_3847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_3858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1020 net1023 VGND VGND VPWR VPWR net1020 sky130_fd_sc_hd__clkbuf_2
Xfanout1031 _05460_ VGND VGND VPWR VPWR net1031 sky130_fd_sc_hd__buf_1
Xfanout1042 _05454_ VGND VGND VPWR VPWR net1042 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1053 _05448_ VGND VGND VPWR VPWR net1053 sky130_fd_sc_hd__buf_1
XFILLER_117_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10168_ net873 net4187 net366 VGND VGND VPWR VPWR _01916_ sky130_fd_sc_hd__mux2_1
XFILLER_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1064 net1065 VGND VGND VPWR VPWR net1064 sky130_fd_sc_hd__clkbuf_2
Xfanout1075 _05438_ VGND VGND VPWR VPWR net1075 sky130_fd_sc_hd__buf_1
Xfanout1086 net1087 VGND VGND VPWR VPWR net1086 sky130_fd_sc_hd__clkbuf_2
Xfanout1097 _05426_ VGND VGND VPWR VPWR net1097 sky130_fd_sc_hd__clkbuf_1
X_10099_ net1792 net728 net642 VGND VGND VPWR VPWR _01848_ sky130_fd_sc_hd__mux2_1
X_13927_ clknet_leaf_39_clk _02556_ VGND VGND VPWR VPWR data_array.data1\[4\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_179_Right_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13858_ clknet_leaf_254_clk _02487_ VGND VGND VPWR VPWR data_array.data1\[3\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12809_ clknet_leaf_32_clk _01503_ VGND VGND VPWR VPWR tag_array.tag1\[0\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_62_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_108_clk clknet_5_27__leaf_clk VGND VGND VPWR VPWR clknet_leaf_108_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_44_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13789_ clknet_leaf_228_clk _02418_ VGND VGND VPWR VPWR data_array.data1\[2\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_06330_ tag_array.tag0\[9\]\[13\] net1608 net1512 tag_array.tag0\[10\]\[13\] VGND
+ VGND VPWR VPWR _03672_ sky130_fd_sc_hd__a22o_1
XFILLER_163_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06261_ net1200 _03603_ _03607_ net1626 VGND VGND VPWR VPWR _03610_ sky130_fd_sc_hd__a22o_1
X_08000_ net1166 _05185_ _05189_ net1214 VGND VGND VPWR VPWR _05191_ sky130_fd_sc_hd__a22o_1
XFILLER_116_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06192_ tag_array.tag0\[12\]\[0\] net1406 net1312 tag_array.tag0\[15\]\[0\] _03546_
+ VGND VGND VPWR VPWR _03547_ sky130_fd_sc_hd__a221o_1
Xhold503 data_array.data0\[0\]\[11\] VGND VGND VPWR VPWR net2154 sky130_fd_sc_hd__dlygate4sd3_1
Xhold514 data_array.data0\[13\]\[49\] VGND VGND VPWR VPWR net2165 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold525 data_array.data1\[8\]\[28\] VGND VGND VPWR VPWR net2176 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold536 data_array.data0\[8\]\[61\] VGND VGND VPWR VPWR net2187 sky130_fd_sc_hd__dlygate4sd3_1
Xhold547 data_array.data0\[2\]\[24\] VGND VGND VPWR VPWR net2198 sky130_fd_sc_hd__dlygate4sd3_1
Xhold558 data_array.data1\[1\]\[42\] VGND VGND VPWR VPWR net2209 sky130_fd_sc_hd__dlygate4sd3_1
X_09951_ net1027 net3744 net372 VGND VGND VPWR VPWR _01700_ sky130_fd_sc_hd__mux2_1
Xhold569 data_array.data0\[1\]\[36\] VGND VGND VPWR VPWR net2220 sky130_fd_sc_hd__dlygate4sd3_1
X_08902_ net896 net2841 net434 VGND VGND VPWR VPWR _00659_ sky130_fd_sc_hd__mux2_1
XFILLER_83_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09882_ net941 net3408 net385 VGND VGND VPWR VPWR _01632_ sky130_fd_sc_hd__mux2_1
XFILLER_170_1022 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08833_ net1767 net913 net447 VGND VGND VPWR VPWR _00591_ sky130_fd_sc_hd__mux2_1
Xhold1203 data_array.data0\[13\]\[15\] VGND VGND VPWR VPWR net2854 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1214 data_array.data1\[9\]\[18\] VGND VGND VPWR VPWR net2865 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1225 tag_array.tag1\[7\]\[22\] VGND VGND VPWR VPWR net2876 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1236 tag_array.tag0\[15\]\[5\] VGND VGND VPWR VPWR net2887 sky130_fd_sc_hd__dlygate4sd3_1
X_08764_ net768 net4534 net450 VGND VGND VPWR VPWR _00523_ sky130_fd_sc_hd__mux2_1
Xhold1247 data_array.data1\[3\]\[31\] VGND VGND VPWR VPWR net2898 sky130_fd_sc_hd__dlygate4sd3_1
X_05976_ data_array.rdata1\[48\] net833 net842 VGND VGND VPWR VPWR _03445_ sky130_fd_sc_hd__a21o_1
Xhold1258 tag_array.tag0\[3\]\[11\] VGND VGND VPWR VPWR net2909 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1269 data_array.data0\[9\]\[16\] VGND VGND VPWR VPWR net2920 sky130_fd_sc_hd__dlygate4sd3_1
X_07715_ _04930_ _04931_ VGND VGND VPWR VPWR _00080_ sky130_fd_sc_hd__or2_1
XFILLER_38_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08695_ net1853 net742 net488 VGND VGND VPWR VPWR _00454_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_140_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07646_ data_array.data1\[0\]\[18\] net1344 net1250 data_array.data1\[3\]\[18\] _04868_
+ VGND VGND VPWR VPWR _04869_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_146_Right_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_101_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07577_ data_array.data1\[13\]\[12\] net1587 net1491 data_array.data1\[14\]\[12\]
+ VGND VGND VPWR VPWR _04806_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_81_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09316_ net714 net2698 net548 VGND VGND VPWR VPWR _01070_ sky130_fd_sc_hd__mux2_1
XFILLER_179_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06528_ tag_array.tag1\[13\]\[6\] net1554 net1458 tag_array.tag1\[14\]\[6\] VGND
+ VGND VPWR VPWR _03852_ sky130_fd_sc_hd__a22o_1
X_09247_ net792 net4608 net573 VGND VGND VPWR VPWR _01001_ sky130_fd_sc_hd__mux2_1
XFILLER_21_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06459_ net1626 _03783_ _03787_ net1201 VGND VGND VPWR VPWR _03790_ sky130_fd_sc_hd__a22o_1
XFILLER_182_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09178_ net768 net2976 net629 VGND VGND VPWR VPWR _00932_ sky130_fd_sc_hd__mux2_1
XFILLER_107_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08129_ data_array.data1\[1\]\[62\] net1605 net1509 data_array.data1\[2\]\[62\] VGND
+ VGND VPWR VPWR _05308_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_79_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11140_ net959 net3649 net549 VGND VGND VPWR VPWR _02883_ sky130_fd_sc_hd__mux2_1
XFILLER_150_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_164_3511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_164_3522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11071_ net2472 net976 net333 VGND VGND VPWR VPWR _02814_ sky130_fd_sc_hd__mux2_1
XFILLER_0_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput101 mem_rdata[11] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_1
Xinput112 mem_rdata[21] VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__clkbuf_1
X_10022_ net999 net3726 net557 VGND VGND VPWR VPWR _01771_ sky130_fd_sc_hd__mux2_1
XFILLER_103_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput123 mem_rdata[31] VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_1
Xinput134 mem_rdata[41] VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_1
XFILLER_49_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput145 mem_rdata[51] VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_1
Xhold2460 tag_array.tag0\[7\]\[4\] VGND VGND VPWR VPWR net4111 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput156 mem_rdata[61] VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__buf_1
Xhold2471 tag_array.tag0\[9\]\[13\] VGND VGND VPWR VPWR net4122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2482 data_array.data0\[15\]\[33\] VGND VGND VPWR VPWR net4133 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2493 data_array.data1\[6\]\[24\] VGND VGND VPWR VPWR net4144 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_5_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1770 data_array.data1\[2\]\[46\] VGND VGND VPWR VPWR net3421 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1781 data_array.data0\[9\]\[36\] VGND VGND VPWR VPWR net3432 sky130_fd_sc_hd__dlygate4sd3_1
X_11973_ clknet_leaf_91_clk _00781_ VGND VGND VPWR VPWR data_array.data0\[4\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1792 data_array.data0\[13\]\[58\] VGND VGND VPWR VPWR net3443 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10924_ net1044 net2558 net528 VGND VGND VPWR VPWR _02669_ sky130_fd_sc_hd__mux2_1
X_13712_ clknet_leaf_19_clk _02341_ VGND VGND VPWR VPWR data_array.data1\[1\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_113_Right_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13643_ clknet_leaf_35_clk _02272_ VGND VGND VPWR VPWR data_array.data1\[15\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_10855_ net1066 net4054 net522 VGND VGND VPWR VPWR _02600_ sky130_fd_sc_hd__mux2_1
XFILLER_112_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13574_ clknet_leaf_33_clk _02203_ VGND VGND VPWR VPWR tag_array.dirty1\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_12_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10786_ net2072 net1086 net502 VGND VGND VPWR VPWR _02531_ sky130_fd_sc_hd__mux2_1
XFILLER_13_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12525_ clknet_leaf_134_clk _01219_ VGND VGND VPWR VPWR tag_array.tag1\[11\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12456_ clknet_leaf_18_clk _01150_ VGND VGND VPWR VPWR data_array.data1\[9\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_136_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_326 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11407_ clknet_leaf_100_clk _00217_ VGND VGND VPWR VPWR tag_array.tag1\[7\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_10_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12387_ clknet_leaf_205_clk _01081_ VGND VGND VPWR VPWR data_array.data0\[14\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_126_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_184_3909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14126_ clknet_leaf_88_clk _02755_ VGND VGND VPWR VPWR data_array.data0\[1\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
X_11338_ net942 net3906 net802 VGND VGND VPWR VPWR _03081_ sky130_fd_sc_hd__mux2_1
XFILLER_107_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14057_ clknet_leaf_74_clk _02686_ VGND VGND VPWR VPWR data_array.data1\[6\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
X_11269_ net952 net4052 net676 VGND VGND VPWR VPWR _03012_ sky130_fd_sc_hd__mux2_1
X_13008_ clknet_leaf_175_clk _01702_ VGND VGND VPWR VPWR data_array.data0\[3\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_37_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05830_ _03338_ _03341_ _03342_ _03346_ VGND VGND VPWR VPWR _03347_ sky130_fd_sc_hd__nor4_1
XFILLER_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05761_ net17 fsm.tag_out1\[17\] VGND VGND VPWR VPWR _03278_ sky130_fd_sc_hd__and2b_1
X_07500_ data_array.data1\[13\]\[5\] net1551 net1455 data_array.data1\[14\]\[5\] VGND
+ VGND VPWR VPWR _04736_ sky130_fd_sc_hd__a22o_1
X_08480_ net813 _05556_ VGND VGND VPWR VPWR _05557_ sky130_fd_sc_hd__and2_4
X_05692_ fsm.tag_out0\[22\] net22 VGND VGND VPWR VPWR _03209_ sky130_fd_sc_hd__and2b_1
X_07431_ data_array.data0\[12\]\[63\] net1357 net1263 data_array.data0\[15\]\[63\]
+ _04672_ VGND VGND VPWR VPWR _04673_ sky130_fd_sc_hd__a221o_1
XFILLER_22_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07362_ net1168 _04605_ _04609_ net1216 VGND VGND VPWR VPWR _04611_ sky130_fd_sc_hd__a22o_1
XFILLER_148_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09101_ net882 net4348 net413 VGND VGND VPWR VPWR _00855_ sky130_fd_sc_hd__mux2_1
XFILLER_31_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06313_ tag_array.tag0\[8\]\[11\] net1402 net1308 tag_array.tag0\[11\]\[11\] _03656_
+ VGND VGND VPWR VPWR _03657_ sky130_fd_sc_hd__a221o_1
XFILLER_176_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07293_ data_array.data0\[1\]\[50\] net1537 net1441 data_array.data0\[2\]\[50\] VGND
+ VGND VPWR VPWR _04548_ sky130_fd_sc_hd__a22o_1
X_09032_ net2125 net896 net418 VGND VGND VPWR VPWR _00787_ sky130_fd_sc_hd__mux2_1
XFILLER_108_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06244_ tag_array.tag0\[5\]\[5\] net1607 net1511 tag_array.tag0\[6\]\[5\] VGND VGND
+ VPWR VPWR _03594_ sky130_fd_sc_hd__a22o_1
Xhold300 data_array.data0\[2\]\[25\] VGND VGND VPWR VPWR net1951 sky130_fd_sc_hd__dlygate4sd3_1
X_06175_ _03530_ _03531_ VGND VGND VPWR VPWR _00181_ sky130_fd_sc_hd__or2_1
Xhold311 data_array.data1\[0\]\[49\] VGND VGND VPWR VPWR net1962 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_11_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold322 data_array.data0\[1\]\[11\] VGND VGND VPWR VPWR net1973 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold333 data_array.data0\[4\]\[44\] VGND VGND VPWR VPWR net1984 sky130_fd_sc_hd__dlygate4sd3_1
Xhold344 data_array.data1\[4\]\[11\] VGND VGND VPWR VPWR net1995 sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 data_array.data0\[8\]\[14\] VGND VGND VPWR VPWR net2006 sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 tag_array.tag1\[8\]\[21\] VGND VGND VPWR VPWR net2017 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold377 data_array.data1\[4\]\[28\] VGND VGND VPWR VPWR net2028 sky130_fd_sc_hd__dlygate4sd3_1
Xhold388 tag_array.dirty1\[8\] VGND VGND VPWR VPWR net2039 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout802 net803 VGND VGND VPWR VPWR net802 sky130_fd_sc_hd__buf_2
Xhold399 data_array.data0\[10\]\[49\] VGND VGND VPWR VPWR net2050 sky130_fd_sc_hd__dlygate4sd3_1
X_09934_ net1092 net4062 net375 VGND VGND VPWR VPWR _01683_ sky130_fd_sc_hd__mux2_1
Xfanout813 net814 VGND VGND VPWR VPWR net813 sky130_fd_sc_hd__buf_2
Xfanout824 net825 VGND VGND VPWR VPWR net824 sky130_fd_sc_hd__clkbuf_2
Xfanout835 net836 VGND VGND VPWR VPWR net835 sky130_fd_sc_hd__buf_12
Xfanout846 net847 VGND VGND VPWR VPWR net846 sky130_fd_sc_hd__buf_6
XFILLER_131_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09865_ net1011 net3566 net378 VGND VGND VPWR VPWR _01615_ sky130_fd_sc_hd__mux2_1
Xfanout857 _05546_ VGND VGND VPWR VPWR net857 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1000 data_array.data0\[5\]\[34\] VGND VGND VPWR VPWR net2651 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout868 net869 VGND VGND VPWR VPWR net868 sky130_fd_sc_hd__clkbuf_2
XFILLER_140_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1011 data_array.data1\[1\]\[33\] VGND VGND VPWR VPWR net2662 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout879 _05536_ VGND VGND VPWR VPWR net879 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1022 data_array.data1\[3\]\[8\] VGND VGND VPWR VPWR net2673 sky130_fd_sc_hd__dlygate4sd3_1
X_08816_ net2001 net983 net442 VGND VGND VPWR VPWR _00574_ sky130_fd_sc_hd__mux2_1
XFILLER_86_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1033 tag_array.tag0\[6\]\[18\] VGND VGND VPWR VPWR net2684 sky130_fd_sc_hd__dlygate4sd3_1
X_09796_ net1026 net3786 net388 VGND VGND VPWR VPWR _01547_ sky130_fd_sc_hd__mux2_1
Xhold1044 tag_array.tag0\[5\]\[10\] VGND VGND VPWR VPWR net2695 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1055 tag_array.tag1\[0\]\[20\] VGND VGND VPWR VPWR net2706 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1066 tag_array.tag0\[15\]\[16\] VGND VGND VPWR VPWR net2717 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1077 data_array.data1\[5\]\[53\] VGND VGND VPWR VPWR net2728 sky130_fd_sc_hd__dlygate4sd3_1
X_08747_ net734 net4099 net455 VGND VGND VPWR VPWR _00506_ sky130_fd_sc_hd__mux2_1
XFILLER_100_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05959_ net135 net1155 _03432_ _03433_ VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__a22o_1
Xhold1088 data_array.data0\[4\]\[0\] VGND VGND VPWR VPWR net2739 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1099 tag_array.tag1\[1\]\[14\] VGND VGND VPWR VPWR net2750 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_53_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08678_ net711 net4293 net492 VGND VGND VPWR VPWR _00437_ sky130_fd_sc_hd__mux2_1
XFILLER_54_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07629_ data_array.data1\[12\]\[17\] net1339 net1245 data_array.data1\[15\]\[17\]
+ _04852_ VGND VGND VPWR VPWR _04853_ sky130_fd_sc_hd__a221o_1
XFILLER_158_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10640_ net2412 net900 net469 VGND VGND VPWR VPWR _02385_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_157_3381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10571_ net922 net4378 net462 VGND VGND VPWR VPWR _02316_ sky130_fd_sc_hd__mux2_1
XFILLER_166_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12310_ clknet_leaf_140_clk _01068_ VGND VGND VPWR VPWR tag_array.tag1\[12\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_13290_ clknet_leaf_224_clk _01920_ VGND VGND VPWR VPWR data_array.data0\[11\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_155_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12241_ clknet_leaf_146_clk _00171_ VGND VGND VPWR VPWR fsm.tag_out1\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_181_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12172_ clknet_leaf_181_clk _00980_ VGND VGND VPWR VPWR tag_array.tag0\[14\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_122_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Left_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11123_ net1024 net3356 net542 VGND VGND VPWR VPWR _02866_ sky130_fd_sc_hd__mux2_1
XFILLER_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11054_ net2464 net1047 net330 VGND VGND VPWR VPWR _02797_ sky130_fd_sc_hd__mux2_1
XFILLER_89_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10005_ net1066 net4040 net561 VGND VGND VPWR VPWR _01754_ sky130_fd_sc_hd__mux2_1
XFILLER_76_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2290 data_array.data1\[14\]\[8\] VGND VGND VPWR VPWR net3941 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_64_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11956_ clknet_leaf_71_clk _00764_ VGND VGND VPWR VPWR data_array.data0\[4\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_177_3757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_177_3768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10907_ net858 net2791 net516 VGND VGND VPWR VPWR _02652_ sky130_fd_sc_hd__mux2_1
X_11887_ clknet_leaf_270_clk _00695_ VGND VGND VPWR VPWR data_array.data0\[5\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10838_ net1832 net878 net506 VGND VGND VPWR VPWR _02583_ sky130_fd_sc_hd__mux2_1
X_13626_ clknet_leaf_3_clk _02255_ VGND VGND VPWR VPWR data_array.data0\[9\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_991 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13557_ clknet_leaf_215_clk _02186_ VGND VGND VPWR VPWR data_array.data1\[0\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
X_10769_ net899 net4460 net490 VGND VGND VPWR VPWR _02514_ sky130_fd_sc_hd__mux2_1
XFILLER_9_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12508_ clknet_leaf_120_clk _01202_ VGND VGND VPWR VPWR data_array.data1\[9\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
X_13488_ clknet_leaf_160_clk _02118_ VGND VGND VPWR VPWR tag_array.tag0\[15\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_173_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12439_ clknet_leaf_234_clk _01133_ VGND VGND VPWR VPWR data_array.data0\[14\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_172_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14109_ clknet_leaf_226_clk _02738_ VGND VGND VPWR VPWR data_array.data0\[1\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_07980_ data_array.data1\[13\]\[49\] net1572 net1476 data_array.data1\[14\]\[49\]
+ VGND VGND VPWR VPWR _05172_ sky130_fd_sc_hd__a22o_1
XFILLER_80_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06931_ data_array.data0\[4\]\[17\] net1339 net1245 data_array.data0\[7\]\[17\] _04218_
+ VGND VGND VPWR VPWR _04219_ sky130_fd_sc_hd__a221o_1
X_09650_ net789 net3651 net612 VGND VGND VPWR VPWR _01402_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06862_ data_array.data0\[13\]\[11\] net1568 net1472 data_array.data0\[14\]\[11\]
+ VGND VGND VPWR VPWR _04156_ sky130_fd_sc_hd__a22o_1
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08601_ net719 net2321 net529 VGND VGND VPWR VPWR _00360_ sky130_fd_sc_hd__mux2_1
X_05813_ _03160_ _03168_ _03190_ fsm.valid0 VGND VGND VPWR VPWR _03330_ sky130_fd_sc_hd__or4b_1
X_09581_ net1026 net3631 net396 VGND VGND VPWR VPWR _01333_ sky130_fd_sc_hd__mux2_1
X_06793_ data_array.data0\[8\]\[5\] net1359 net1265 data_array.data0\[11\]\[5\] _04092_
+ VGND VGND VPWR VPWR _04093_ sky130_fd_sc_hd__a221o_1
X_08532_ net1463 net1200 net814 net1702 VGND VGND VPWR VPWR _00305_ sky130_fd_sc_hd__a31o_1
X_05744_ net24 fsm.tag_out1\[23\] VGND VGND VPWR VPWR _03261_ sky130_fd_sc_hd__and2b_1
XFILLER_24_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08463_ net158 net93 net1644 VGND VGND VPWR VPWR _05545_ sky130_fd_sc_hd__mux2_1
XFILLER_91_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05675_ _03181_ _03186_ _03191_ VGND VGND VPWR VPWR _03192_ sky130_fd_sc_hd__or3_1
XFILLER_23_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07414_ data_array.data0\[5\]\[61\] net1548 net1452 data_array.data0\[6\]\[61\] VGND
+ VGND VPWR VPWR _04658_ sky130_fd_sc_hd__a22o_1
X_08394_ net133 net68 net1648 VGND VGND VPWR VPWR _05499_ sky130_fd_sc_hd__mux2_1
XFILLER_51_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07345_ data_array.data0\[0\]\[55\] net1343 net1249 data_array.data0\[3\]\[55\] _04594_
+ VGND VGND VPWR VPWR _04595_ sky130_fd_sc_hd__a221o_1
XFILLER_149_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_30_clk clknet_5_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_30_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_98_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07276_ data_array.data0\[13\]\[49\] net1571 net1475 data_array.data0\[14\]\[49\]
+ VGND VGND VPWR VPWR _04532_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_59_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09015_ net1896 net964 net424 VGND VGND VPWR VPWR _00770_ sky130_fd_sc_hd__mux2_1
X_06227_ tag_array.tag0\[4\]\[3\] net1371 net1277 tag_array.tag0\[7\]\[3\] _03578_
+ VGND VGND VPWR VPWR _03579_ sky130_fd_sc_hd__a221o_1
XFILLER_163_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold130 data_array.data1\[4\]\[13\] VGND VGND VPWR VPWR net1781 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold141 tag_array.tag1\[8\]\[16\] VGND VGND VPWR VPWR net1792 sky130_fd_sc_hd__dlygate4sd3_1
X_06158_ net26 net27 VGND VGND VPWR VPWR _03515_ sky130_fd_sc_hd__and2_2
XFILLER_104_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold152 data_array.data0\[4\]\[19\] VGND VGND VPWR VPWR net1803 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 data_array.data0\[2\]\[35\] VGND VGND VPWR VPWR net1814 sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 data_array.data0\[0\]\[21\] VGND VGND VPWR VPWR net1825 sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 data_array.data0\[8\]\[62\] VGND VGND VPWR VPWR net1836 sky130_fd_sc_hd__dlygate4sd3_1
X_06089_ data_array.rdata0\[4\] net1139 net1115 data_array.rdata1\[4\] VGND VGND VPWR
+ VPWR net307 sky130_fd_sc_hd__a22o_1
Xhold196 data_array.data1\[1\]\[50\] VGND VGND VPWR VPWR net1847 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout610 net611 VGND VGND VPWR VPWR net610 sky130_fd_sc_hd__buf_4
Xfanout1608 net1609 VGND VGND VPWR VPWR net1608 sky130_fd_sc_hd__clkbuf_4
Xfanout621 _05567_ VGND VGND VPWR VPWR net621 sky130_fd_sc_hd__buf_4
XFILLER_132_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1619 net1620 VGND VGND VPWR VPWR net1619 sky130_fd_sc_hd__buf_4
Xfanout632 _05560_ VGND VGND VPWR VPWR net632 sky130_fd_sc_hd__buf_4
X_09917_ net738 net3853 net603 VGND VGND VPWR VPWR _01667_ sky130_fd_sc_hd__mux2_1
Xfanout643 net644 VGND VGND VPWR VPWR net643 sky130_fd_sc_hd__clkbuf_4
Xfanout654 _05551_ VGND VGND VPWR VPWR net654 sky130_fd_sc_hd__buf_4
Xfanout665 net666 VGND VGND VPWR VPWR net665 sky130_fd_sc_hd__clkbuf_8
Xclkbuf_leaf_97_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_97_clk sky130_fd_sc_hd__clkbuf_8
Xfanout676 _05548_ VGND VGND VPWR VPWR net676 sky130_fd_sc_hd__buf_4
XFILLER_19_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout687 net690 VGND VGND VPWR VPWR net687 sky130_fd_sc_hd__buf_4
X_09848_ net1077 net2992 net379 VGND VGND VPWR VPWR _01598_ sky130_fd_sc_hd__mux2_1
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout698 net699 VGND VGND VPWR VPWR net698 sky130_fd_sc_hd__clkbuf_2
XFILLER_100_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_996 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09779_ net1092 net3492 net391 VGND VGND VPWR VPWR _01530_ sky130_fd_sc_hd__mux2_1
XFILLER_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11810_ clknet_leaf_94_clk _00618_ VGND VGND VPWR VPWR data_array.data0\[7\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_159_3410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ clknet_leaf_138_clk _01484_ VGND VGND VPWR VPWR tag_array.tag1\[10\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_163_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_159_3421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11741_ clknet_leaf_86_clk _00549_ VGND VGND VPWR VPWR data_array.data0\[8\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11672_ clknet_leaf_133_clk _00480_ VGND VGND VPWR VPWR tag_array.tag1\[1\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_14460_ clknet_leaf_78_clk _03083_ VGND VGND VPWR VPWR data_array.data1\[7\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10623_ net1861 net968 net468 VGND VGND VPWR VPWR _02368_ sky130_fd_sc_hd__mux2_1
X_13411_ clknet_leaf_37_clk _02041_ VGND VGND VPWR VPWR data_array.data1\[8\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_14391_ clknet_leaf_260_clk _03014_ VGND VGND VPWR VPWR data_array.data1\[10\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_12_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_172_3665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_21_clk clknet_5_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_8
X_13342_ clknet_leaf_3_clk _01972_ VGND VGND VPWR VPWR data_array.data0\[10\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10554_ net991 net3075 net461 VGND VGND VPWR VPWR _02299_ sky130_fd_sc_hd__mux2_1
XFILLER_6_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_133_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_656 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13273_ clknet_leaf_23_clk _01903_ VGND VGND VPWR VPWR data_array.data0\[11\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
X_10485_ net1006 net2734 net345 VGND VGND VPWR VPWR _02230_ sky130_fd_sc_hd__mux2_1
X_12224_ clknet_leaf_183_clk _00177_ VGND VGND VPWR VPWR fsm.tag_out1\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12155_ clknet_leaf_154_clk _00963_ VGND VGND VPWR VPWR tag_array.tag0\[13\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_151_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11106_ net1095 net2984 net549 VGND VGND VPWR VPWR _02849_ sky130_fd_sc_hd__mux2_1
X_12086_ clknet_leaf_264_clk _00894_ VGND VGND VPWR VPWR data_array.data1\[14\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_34_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_88_clk clknet_5_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_88_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_34_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11037_ _05352_ net807 VGND VGND VPWR VPWR _03133_ sky130_fd_sc_hd__and2_4
XFILLER_49_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_179_3808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12988_ clknet_leaf_48_clk _01682_ VGND VGND VPWR VPWR data_array.data0\[3\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_11939_ clknet_leaf_206_clk _00747_ VGND VGND VPWR VPWR data_array.data0\[4\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_928 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13609_ clknet_leaf_11_clk _02238_ VGND VGND VPWR VPWR data_array.data0\[9\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_12_clk clknet_5_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_8
X_07130_ net1193 _04393_ _04397_ net1619 VGND VGND VPWR VPWR _04400_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_31_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07061_ data_array.data0\[8\]\[29\] net1379 net1285 data_array.data0\[11\]\[29\]
+ _04336_ VGND VGND VPWR VPWR _04337_ sky130_fd_sc_hd__a221o_1
XFILLER_145_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06012_ data_array.rdata1\[60\] net1657 net843 VGND VGND VPWR VPWR _03469_ sky130_fd_sc_hd__a21o_1
Xoutput202 net202 VGND VGND VPWR VPWR cpu_rdata[43] sky130_fd_sc_hd__clkbuf_4
Xoutput213 net213 VGND VGND VPWR VPWR cpu_rdata[53] sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_93_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput224 net224 VGND VGND VPWR VPWR cpu_rdata[63] sky130_fd_sc_hd__buf_2
Xoutput235 net235 VGND VGND VPWR VPWR mem_addr[14] sky130_fd_sc_hd__buf_2
XFILLER_142_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput246 net246 VGND VGND VPWR VPWR mem_addr[24] sky130_fd_sc_hd__buf_2
Xoutput257 net257 VGND VGND VPWR VPWR mem_addr[5] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput268 net268 VGND VGND VPWR VPWR mem_wdata[14] sky130_fd_sc_hd__buf_2
Xoutput279 net279 VGND VGND VPWR VPWR mem_wdata[24] sky130_fd_sc_hd__buf_2
XFILLER_141_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07963_ data_array.data1\[12\]\[47\] net1397 net1303 data_array.data1\[15\]\[47\]
+ _05156_ VGND VGND VPWR VPWR _05157_ sky130_fd_sc_hd__a221o_1
XFILLER_141_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_71_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_79_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_79_clk sky130_fd_sc_hd__clkbuf_8
X_06914_ data_array.data0\[8\]\[16\] net1357 net1263 data_array.data0\[11\]\[16\]
+ _04202_ VGND VGND VPWR VPWR _04203_ sky130_fd_sc_hd__a221o_1
X_09702_ net780 net2526 net609 VGND VGND VPWR VPWR _01454_ sky130_fd_sc_hd__mux2_1
X_07894_ data_array.data1\[5\]\[41\] net1525 net1429 data_array.data1\[6\]\[41\] VGND
+ VGND VPWR VPWR _05094_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_74_Left_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09633_ net755 net3805 net616 VGND VGND VPWR VPWR _01385_ sky130_fd_sc_hd__mux2_1
X_06845_ net1178 _04135_ _04139_ net1226 VGND VGND VPWR VPWR _04141_ sky130_fd_sc_hd__a22o_1
XFILLER_83_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09564_ net1092 net4301 net399 VGND VGND VPWR VPWR _01316_ sky130_fd_sc_hd__mux2_1
X_06776_ data_array.data0\[1\]\[3\] net1567 net1471 data_array.data0\[2\]\[3\] VGND
+ VGND VPWR VPWR _04078_ sky130_fd_sc_hd__a22o_1
X_08515_ _03514_ _03527_ net823 VGND VGND VPWR VPWR _05581_ sky130_fd_sc_hd__or3_1
X_05727_ fsm.valid1 _03242_ _03243_ VGND VGND VPWR VPWR _03244_ sky130_fd_sc_hd__and3_1
X_09495_ net748 net3536 net625 VGND VGND VPWR VPWR _01248_ sky130_fd_sc_hd__mux2_1
XFILLER_169_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08446_ net1125 _05533_ VGND VGND VPWR VPWR _05534_ sky130_fd_sc_hd__and2_1
X_05658_ fsm.tag_out0\[19\] net19 VGND VGND VPWR VPWR _03175_ sky130_fd_sc_hd__and2b_1
XFILLER_24_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08377_ net1124 _05487_ VGND VGND VPWR VPWR _05488_ sky130_fd_sc_hd__and2_1
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07328_ net1615 _04573_ _04577_ net1189 VGND VGND VPWR VPWR _04580_ sky130_fd_sc_hd__a22o_1
XFILLER_177_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_83_Left_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07259_ data_array.data0\[12\]\[47\] net1387 net1293 data_array.data0\[15\]\[47\]
+ _04516_ VGND VGND VPWR VPWR _04517_ sky130_fd_sc_hd__a221o_1
XFILLER_180_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10270_ net1980 net1082 net641 VGND VGND VPWR VPWR _02017_ sky130_fd_sc_hd__mux2_1
XFILLER_105_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1405 net1406 VGND VGND VPWR VPWR net1405 sky130_fd_sc_hd__clkbuf_4
Xfanout1416 net1422 VGND VGND VPWR VPWR net1416 sky130_fd_sc_hd__buf_2
Xfanout1427 net1428 VGND VGND VPWR VPWR net1427 sky130_fd_sc_hd__clkbuf_4
Xfanout440 net441 VGND VGND VPWR VPWR net440 sky130_fd_sc_hd__buf_4
XFILLER_63_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1438 net1440 VGND VGND VPWR VPWR net1438 sky130_fd_sc_hd__clkbuf_4
Xfanout1449 net1450 VGND VGND VPWR VPWR net1449 sky130_fd_sc_hd__clkbuf_4
Xfanout451 _05606_ VGND VGND VPWR VPWR net451 sky130_fd_sc_hd__buf_4
Xfanout462 net465 VGND VGND VPWR VPWR net462 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_92_Left_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13960_ clknet_leaf_227_clk _02589_ VGND VGND VPWR VPWR data_array.data1\[5\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout473 net474 VGND VGND VPWR VPWR net473 sky130_fd_sc_hd__buf_2
XFILLER_24_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout484 net486 VGND VGND VPWR VPWR net484 sky130_fd_sc_hd__clkbuf_8
XFILLER_171_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout495 _05601_ VGND VGND VPWR VPWR net495 sky130_fd_sc_hd__clkbuf_4
XFILLER_47_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12911_ clknet_leaf_63_clk _01605_ VGND VGND VPWR VPWR data_array.data0\[13\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13891_ clknet_leaf_41_clk _02520_ VGND VGND VPWR VPWR data_array.data1\[3\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12842_ clknet_leaf_111_clk _01536_ VGND VGND VPWR VPWR data_array.data0\[12\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_174_3705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ clknet_leaf_157_clk _01467_ VGND VGND VPWR VPWR tag_array.tag0\[6\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11724_ clknet_leaf_162_clk _00532_ VGND VGND VPWR VPWR tag_array.tag0\[9\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_14443_ clknet_leaf_220_clk _03066_ VGND VGND VPWR VPWR data_array.data1\[7\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_80_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11655_ clknet_leaf_100_clk _00463_ VGND VGND VPWR VPWR tag_array.tag1\[2\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_80_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10606_ net1862 net1038 net471 VGND VGND VPWR VPWR _02351_ sky130_fd_sc_hd__mux2_1
X_11586_ clknet_leaf_233_clk _00394_ VGND VGND VPWR VPWR tag_array.tag1\[4\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14374_ clknet_leaf_89_clk _02997_ VGND VGND VPWR VPWR data_array.data1\[10\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_167_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10537_ net1056 net2090 net457 VGND VGND VPWR VPWR _02282_ sky130_fd_sc_hd__mux2_1
X_13325_ clknet_leaf_10_clk _01955_ VGND VGND VPWR VPWR data_array.data0\[10\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_155_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13256_ clknet_leaf_54_clk _01886_ VGND VGND VPWR VPWR data_array.data0\[11\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_10468_ net1073 net3471 net348 VGND VGND VPWR VPWR _02213_ sky130_fd_sc_hd__mux2_1
X_12207_ clknet_leaf_182_clk _00136_ VGND VGND VPWR VPWR fsm.tag_out0\[14\] sky130_fd_sc_hd__dfxtp_1
X_13187_ clknet_leaf_80_clk _00080_ VGND VGND VPWR VPWR data_array.rdata1\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_9_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10399_ net1766 net1056 net664 VGND VGND VPWR VPWR _02145_ sky130_fd_sc_hd__mux2_1
X_12138_ clknet_leaf_171_clk _00946_ VGND VGND VPWR VPWR tag_array.tag0\[12\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_96_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12069_ clknet_leaf_59_clk _00877_ VGND VGND VPWR VPWR data_array.data1\[14\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_1_clk clknet_5_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_38_836 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06630_ tag_array.tag1\[0\]\[15\] net1385 net1291 tag_array.tag1\[3\]\[15\] _03944_
+ VGND VGND VPWR VPWR _03945_ sky130_fd_sc_hd__a221o_1
XFILLER_37_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06561_ tag_array.tag1\[9\]\[9\] net1609 net1513 tag_array.tag1\[10\]\[9\] VGND VGND
+ VPWR VPWR _03882_ sky130_fd_sc_hd__a22o_1
X_08300_ net1925 net1076 net687 VGND VGND VPWR VPWR _00229_ sky130_fd_sc_hd__mux2_1
X_09280_ net761 net4037 net565 VGND VGND VPWR VPWR _01034_ sky130_fd_sc_hd__mux2_1
X_06492_ net1619 _03813_ _03817_ net1193 VGND VGND VPWR VPWR _03820_ sky130_fd_sc_hd__a22o_1
XFILLER_33_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08231_ fsm.tag_out1\[12\] _05359_ _05364_ fsm.tag_out0\[12\] _05388_ VGND VGND VPWR
+ VPWR _05389_ sky130_fd_sc_hd__a221o_2
XTAP_TAPCELL_ROW_95_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08162_ tag_array.dirty0\[5\] net1593 net1497 tag_array.dirty0\[6\] VGND VGND VPWR
+ VPWR _05338_ sky130_fd_sc_hd__a22o_1
XFILLER_146_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07113_ data_array.data0\[5\]\[34\] net1531 net1435 data_array.data0\[6\]\[34\] VGND
+ VGND VPWR VPWR _04384_ sky130_fd_sc_hd__a22o_1
XFILLER_147_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08093_ data_array.data1\[0\]\[59\] net1381 net1287 data_array.data1\[3\]\[59\] _05274_
+ VGND VGND VPWR VPWR _05275_ sky130_fd_sc_hd__a221o_1
XFILLER_134_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload50 clknet_leaf_246_clk VGND VGND VPWR VPWR clkload50/X sky130_fd_sc_hd__clkbuf_4
XFILLER_118_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07044_ _04320_ _04321_ VGND VGND VPWR VPWR _00019_ sky130_fd_sc_hd__or2_1
Xclkload61 clknet_leaf_27_clk VGND VGND VPWR VPWR clkload61/Y sky130_fd_sc_hd__inv_8
XFILLER_134_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload72 clknet_leaf_238_clk VGND VGND VPWR VPWR clkload72/Y sky130_fd_sc_hd__inv_8
XFILLER_127_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload83 clknet_leaf_43_clk VGND VGND VPWR VPWR clkload83/Y sky130_fd_sc_hd__inv_6
XFILLER_161_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload94 clknet_leaf_56_clk VGND VGND VPWR VPWR clkload94/Y sky130_fd_sc_hd__inv_6
XFILLER_86_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2801 data_array.data0\[3\]\[51\] VGND VGND VPWR VPWR net4452 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2812 data_array.data0\[14\]\[53\] VGND VGND VPWR VPWR net4463 sky130_fd_sc_hd__dlygate4sd3_1
X_08995_ net1939 net1047 net420 VGND VGND VPWR VPWR _00750_ sky130_fd_sc_hd__mux2_1
Xhold2823 data_array.data1\[7\]\[25\] VGND VGND VPWR VPWR net4474 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2834 tag_array.tag0\[10\]\[4\] VGND VGND VPWR VPWR net4485 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2845 tag_array.tag0\[9\]\[3\] VGND VGND VPWR VPWR net4496 sky130_fd_sc_hd__dlygate4sd3_1
X_07946_ _05140_ _05141_ VGND VGND VPWR VPWR _00103_ sky130_fd_sc_hd__or2_1
XFILLER_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2856 tag_array.tag0\[5\]\[5\] VGND VGND VPWR VPWR net4507 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2867 data_array.data1\[11\]\[29\] VGND VGND VPWR VPWR net4518 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2878 tag_array.tag1\[5\]\[13\] VGND VGND VPWR VPWR net4529 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2889 tag_array.tag0\[11\]\[19\] VGND VGND VPWR VPWR net4540 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07877_ data_array.data1\[4\]\[39\] net1347 net1253 data_array.data1\[7\]\[39\] _05078_
+ VGND VGND VPWR VPWR _05079_ sky130_fd_sc_hd__a221o_1
XFILLER_56_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09616_ net885 net2951 net395 VGND VGND VPWR VPWR _01368_ sky130_fd_sc_hd__mux2_1
X_06828_ data_array.data0\[4\]\[8\] net1345 net1251 data_array.data0\[7\]\[8\] _04124_
+ VGND VGND VPWR VPWR _04125_ sky130_fd_sc_hd__a221o_1
XFILLER_56_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06759_ data_array.data0\[13\]\[2\] net1528 net1432 data_array.data0\[14\]\[2\] VGND
+ VGND VPWR VPWR _04062_ sky130_fd_sc_hd__a22o_1
XFILLER_93_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_104_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09547_ net739 net4227 net620 VGND VGND VPWR VPWR _01300_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09478_ net715 net4465 net655 VGND VGND VPWR VPWR _01231_ sky130_fd_sc_hd__mux2_1
XFILLER_180_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_568 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08429_ net1949 net904 net686 VGND VGND VPWR VPWR _00272_ sky130_fd_sc_hd__mux2_1
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload0 clknet_5_0__leaf_clk VGND VGND VPWR VPWR clkload0/X sky130_fd_sc_hd__clkbuf_8
X_11440_ clknet_leaf_53_clk _00250_ VGND VGND VPWR VPWR data_array.data0\[0\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_126_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_966 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11371_ net1646 net2901 net622 VGND VGND VPWR VPWR _03114_ sky130_fd_sc_hd__mux2_1
XFILLER_138_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13110_ clknet_leaf_203_clk _01804_ VGND VGND VPWR VPWR data_array.data1\[13\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
X_10322_ net1954 net874 net639 VGND VGND VPWR VPWR _02069_ sky130_fd_sc_hd__mux2_1
XFILLER_30_1071 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14090_ clknet_leaf_247_clk _02719_ VGND VGND VPWR VPWR data_array.data0\[1\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_124_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13041_ clknet_leaf_12_clk _01735_ VGND VGND VPWR VPWR data_array.data0\[3\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
X_10253_ net732 net3149 net595 VGND VGND VPWR VPWR _02000_ sky130_fd_sc_hd__mux2_1
Xclkbuf_5_29__f_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_5_29__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_167_3564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_3575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1202 net1203 VGND VGND VPWR VPWR net1202 sky130_fd_sc_hd__buf_4
XFILLER_132_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10184_ net1069 net3087 net360 VGND VGND VPWR VPWR _01931_ sky130_fd_sc_hd__mux2_1
Xfanout1213 net1215 VGND VGND VPWR VPWR net1213 sky130_fd_sc_hd__buf_4
XFILLER_182_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1224 net1225 VGND VGND VPWR VPWR net1224 sky130_fd_sc_hd__buf_4
Xfanout1235 net1237 VGND VGND VPWR VPWR net1235 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_128_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1246 net1248 VGND VGND VPWR VPWR net1246 sky130_fd_sc_hd__clkbuf_4
XFILLER_94_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1257 net1258 VGND VGND VPWR VPWR net1257 sky130_fd_sc_hd__clkbuf_2
Xfanout1268 net1269 VGND VGND VPWR VPWR net1268 sky130_fd_sc_hd__clkbuf_4
Xfanout1279 net1280 VGND VGND VPWR VPWR net1279 sky130_fd_sc_hd__clkbuf_4
X_13943_ clknet_leaf_78_clk _02572_ VGND VGND VPWR VPWR data_array.data1\[4\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13874_ clknet_leaf_88_clk _02503_ VGND VGND VPWR VPWR data_array.data1\[3\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12825_ clknet_leaf_187_clk _01519_ VGND VGND VPWR VPWR tag_array.tag1\[0\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_12756_ clknet_leaf_186_clk _01450_ VGND VGND VPWR VPWR tag_array.tag0\[5\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_11707_ clknet_leaf_130_clk _00515_ VGND VGND VPWR VPWR tag_array.tag1\[15\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_12687_ clknet_leaf_146_clk _01381_ VGND VGND VPWR VPWR tag_array.tag0\[8\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_147_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14426_ clknet_leaf_116_clk _03049_ VGND VGND VPWR VPWR data_array.data1\[7\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_11638_ clknet_leaf_193_clk _00446_ VGND VGND VPWR VPWR tag_array.tag1\[2\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_42_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14357_ clknet_leaf_81_clk _02980_ VGND VGND VPWR VPWR data_array.data1\[10\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_11569_ clknet_leaf_103_clk _00377_ VGND VGND VPWR VPWR tag_array.tag1\[5\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold707 tag_array.tag0\[10\]\[20\] VGND VGND VPWR VPWR net2358 sky130_fd_sc_hd__dlygate4sd3_1
X_13308_ clknet_leaf_246_clk _01938_ VGND VGND VPWR VPWR data_array.data0\[10\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold718 tag_array.tag0\[14\]\[24\] VGND VGND VPWR VPWR net2369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold729 data_array.data1\[8\]\[44\] VGND VGND VPWR VPWR net2380 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14288_ clknet_leaf_19_clk _02917_ VGND VGND VPWR VPWR data_array.data1\[11\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_90_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_139_Left_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13239_ clknet_leaf_104_clk _01869_ VGND VGND VPWR VPWR data_array.data0\[11\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_170_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2108 tag_array.tag0\[5\]\[2\] VGND VGND VPWR VPWR net3759 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_124_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2119 data_array.data1\[12\]\[0\] VGND VGND VPWR VPWR net3770 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07800_ data_array.data1\[4\]\[32\] net1330 net1236 data_array.data1\[7\]\[32\] _05008_
+ VGND VGND VPWR VPWR _05009_ sky130_fd_sc_hd__a221o_1
X_08780_ net704 net2503 net450 VGND VGND VPWR VPWR _00539_ sky130_fd_sc_hd__mux2_1
XFILLER_85_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1407 tag_array.tag0\[11\]\[17\] VGND VGND VPWR VPWR net3058 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1418 data_array.data1\[11\]\[7\] VGND VGND VPWR VPWR net3069 sky130_fd_sc_hd__dlygate4sd3_1
X_05992_ net147 net1150 _03454_ _03455_ VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__a22o_1
XFILLER_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_127_Right_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1429 tag_array.tag1\[8\]\[19\] VGND VGND VPWR VPWR net3080 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07731_ data_array.data1\[13\]\[26\] net1525 net1429 data_array.data1\[14\]\[26\]
+ VGND VGND VPWR VPWR _04946_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_88_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_88_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07662_ data_array.data1\[12\]\[20\] net1419 net1325 data_array.data1\[15\]\[20\]
+ _04882_ VGND VGND VPWR VPWR _04883_ sky130_fd_sc_hd__a221o_1
XFILLER_77_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06613_ net1210 _03923_ _03927_ net1636 VGND VGND VPWR VPWR _03930_ sky130_fd_sc_hd__a22o_1
X_09401_ net1063 net3158 net587 VGND VGND VPWR VPWR _01154_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_148_Left_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07593_ net1219 _04815_ _04819_ net1171 VGND VGND VPWR VPWR _04821_ sky130_fd_sc_hd__a22o_1
XFILLER_53_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06544_ tag_array.tag1\[12\]\[7\] net1420 net1326 tag_array.tag1\[15\]\[7\] _03866_
+ VGND VGND VPWR VPWR _03867_ sky130_fd_sc_hd__a221o_1
X_09332_ net1072 net2589 net407 VGND VGND VPWR VPWR _01085_ sky130_fd_sc_hd__mux2_1
XFILLER_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09263_ net729 net3335 net576 VGND VGND VPWR VPWR _01017_ sky130_fd_sc_hd__mux2_1
X_06475_ tag_array.tag1\[5\]\[1\] net1575 net1479 tag_array.tag1\[6\]\[1\] VGND VGND
+ VPWR VPWR _03804_ sky130_fd_sc_hd__a22o_1
X_08214_ net766 net3327 net806 VGND VGND VPWR VPWR _00202_ sky130_fd_sc_hd__mux2_1
X_09194_ net705 net3289 net629 VGND VGND VPWR VPWR _00948_ sky130_fd_sc_hd__mux2_1
X_08145_ tag_array.dirty1\[13\] net1574 net1478 tag_array.dirty1\[14\] VGND VGND VPWR
+ VPWR _05322_ sky130_fd_sc_hd__a22o_1
XFILLER_146_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_157_Left_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08076_ net1190 _05253_ _05257_ net1617 VGND VGND VPWR VPWR _05260_ sky130_fd_sc_hd__a22o_1
Xclkload150 clknet_leaf_227_clk VGND VGND VPWR VPWR clkload150/Y sky130_fd_sc_hd__inv_6
XFILLER_107_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload161 clknet_leaf_174_clk VGND VGND VPWR VPWR clkload161/Y sky130_fd_sc_hd__bufinv_16
Xclkload172 clknet_leaf_197_clk VGND VGND VPWR VPWR clkload172/Y sky130_fd_sc_hd__inv_6
XFILLER_20_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07027_ data_array.data0\[13\]\[26\] net1527 net1431 data_array.data0\[14\]\[26\]
+ VGND VGND VPWR VPWR _04306_ sky130_fd_sc_hd__a22o_1
Xclkload183 clknet_leaf_184_clk VGND VGND VPWR VPWR clkload183/Y sky130_fd_sc_hd__clkinv_4
Xclkload194 clknet_leaf_103_clk VGND VGND VPWR VPWR clkload194/Y sky130_fd_sc_hd__bufinv_16
XFILLER_162_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_927 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2620 data_array.data0\[10\]\[6\] VGND VGND VPWR VPWR net4271 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2631 tag_array.dirty1\[10\] VGND VGND VPWR VPWR net4282 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_145_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2642 tag_array.tag1\[3\]\[20\] VGND VGND VPWR VPWR net4293 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2653 data_array.data1\[3\]\[52\] VGND VGND VPWR VPWR net4304 sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ net807 _05580_ VGND VGND VPWR VPWR _05610_ sky130_fd_sc_hd__and2_1
Xhold45 tag_array.valid1\[3\] VGND VGND VPWR VPWR net1696 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold56 tag_array.valid1\[13\] VGND VGND VPWR VPWR net1707 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2664 data_array.data0\[11\]\[7\] VGND VGND VPWR VPWR net4315 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2675 data_array.data1\[14\]\[6\] VGND VGND VPWR VPWR net4326 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold67 tag_array.valid0\[12\] VGND VGND VPWR VPWR net1718 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1930 tag_array.tag0\[12\]\[0\] VGND VGND VPWR VPWR net3581 sky130_fd_sc_hd__dlygate4sd3_1
X_07929_ data_array.data1\[13\]\[44\] net1589 net1493 data_array.data1\[14\]\[44\]
+ VGND VGND VPWR VPWR _05126_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_162_3472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold78 data_array.data0\[0\]\[17\] VGND VGND VPWR VPWR net1729 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1941 tag_array.tag1\[6\]\[6\] VGND VGND VPWR VPWR net3592 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2686 tag_array.tag0\[1\]\[7\] VGND VGND VPWR VPWR net4337 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_162_3483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2697 data_array.data0\[6\]\[57\] VGND VGND VPWR VPWR net4348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1952 tag_array.tag1\[15\]\[11\] VGND VGND VPWR VPWR net3603 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold89 data_array.data0\[8\]\[19\] VGND VGND VPWR VPWR net1740 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1963 data_array.data0\[11\]\[43\] VGND VGND VPWR VPWR net3614 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_166_Left_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1974 tag_array.tag1\[8\]\[15\] VGND VGND VPWR VPWR net3625 sky130_fd_sc_hd__dlygate4sd3_1
X_10940_ net980 net4487 net526 VGND VGND VPWR VPWR _02685_ sky130_fd_sc_hd__mux2_1
Xhold1985 data_array.data1\[13\]\[53\] VGND VGND VPWR VPWR net3636 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1996 data_array.data0\[3\]\[26\] VGND VGND VPWR VPWR net3647 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_123_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10871_ net1000 net3355 net516 VGND VGND VPWR VPWR _02616_ sky130_fd_sc_hd__mux2_1
X_12610_ clknet_leaf_108_clk _01304_ VGND VGND VPWR VPWR tag_array.tag0\[0\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_13590_ clknet_leaf_64_clk _02219_ VGND VGND VPWR VPWR data_array.data0\[9\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12541_ clknet_leaf_130_clk _01235_ VGND VGND VPWR VPWR tag_array.tag1\[11\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_101_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12472_ clknet_leaf_89_clk _01166_ VGND VGND VPWR VPWR data_array.data1\[9\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_175_Left_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14211_ clknet_leaf_52_clk _02840_ VGND VGND VPWR VPWR data_array.data0\[2\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
X_11423_ clknet_leaf_94_clk _00233_ VGND VGND VPWR VPWR data_array.data0\[0\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_169_3604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_169_3615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_9 _00158_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11354_ net878 net3556 net799 VGND VGND VPWR VPWR _03097_ sky130_fd_sc_hd__mux2_1
X_14142_ clknet_leaf_221_clk _02771_ VGND VGND VPWR VPWR data_array.data0\[1\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_180_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10305_ net2239 net942 net641 VGND VGND VPWR VPWR _02052_ sky130_fd_sc_hd__mux2_1
XFILLER_4_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11285_ net891 net3406 net675 VGND VGND VPWR VPWR _03028_ sky130_fd_sc_hd__mux2_1
X_14073_ clknet_leaf_55_clk _02702_ VGND VGND VPWR VPWR data_array.data1\[6\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
X_10236_ net861 net2122 net361 VGND VGND VPWR VPWR _01983_ sky130_fd_sc_hd__mux2_1
X_13024_ clknet_leaf_235_clk _01718_ VGND VGND VPWR VPWR data_array.data0\[3\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout1010 net1011 VGND VGND VPWR VPWR net1010 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_182_3848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1021 net1022 VGND VGND VPWR VPWR net1021 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_182_3859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1032 net1033 VGND VGND VPWR VPWR net1032 sky130_fd_sc_hd__clkbuf_2
X_10167_ net876 net4220 net365 VGND VGND VPWR VPWR _01915_ sky130_fd_sc_hd__mux2_1
Xfanout1043 _05454_ VGND VGND VPWR VPWR net1043 sky130_fd_sc_hd__buf_1
Xfanout1054 _05448_ VGND VGND VPWR VPWR net1054 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1065 _05442_ VGND VGND VPWR VPWR net1065 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1076 _05436_ VGND VGND VPWR VPWR net1076 sky130_fd_sc_hd__clkbuf_2
Xfanout1087 _05432_ VGND VGND VPWR VPWR net1087 sky130_fd_sc_hd__dlymetal6s2s_1
X_10098_ net3625 net731 net639 VGND VGND VPWR VPWR _01847_ sky130_fd_sc_hd__mux2_1
XFILLER_47_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1098 net1099 VGND VGND VPWR VPWR net1098 sky130_fd_sc_hd__clkbuf_2
XFILLER_48_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13926_ clknet_leaf_69_clk _02555_ VGND VGND VPWR VPWR data_array.data1\[4\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13857_ clknet_leaf_267_clk _02486_ VGND VGND VPWR VPWR data_array.data1\[3\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12808_ clknet_leaf_99_clk _01502_ VGND VGND VPWR VPWR tag_array.tag1\[0\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_13788_ clknet_leaf_122_clk _02417_ VGND VGND VPWR VPWR data_array.data1\[2\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_44_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12739_ clknet_leaf_143_clk _01433_ VGND VGND VPWR VPWR tag_array.tag0\[5\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06260_ tag_array.tag0\[0\]\[6\] net1373 net1280 tag_array.tag0\[3\]\[6\] _03608_
+ VGND VGND VPWR VPWR _03609_ sky130_fd_sc_hd__a221o_1
XFILLER_176_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14409_ clknet_leaf_41_clk _03032_ VGND VGND VPWR VPWR data_array.data1\[10\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
X_06191_ tag_array.tag0\[13\]\[0\] net1596 net1500 tag_array.tag0\[14\]\[0\] VGND
+ VGND VPWR VPWR _03546_ sky130_fd_sc_hd__a22o_1
XFILLER_128_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold504 data_array.data1\[8\]\[31\] VGND VGND VPWR VPWR net2155 sky130_fd_sc_hd__dlygate4sd3_1
Xhold515 data_array.data1\[2\]\[17\] VGND VGND VPWR VPWR net2166 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold526 data_array.data1\[0\]\[32\] VGND VGND VPWR VPWR net2177 sky130_fd_sc_hd__dlygate4sd3_1
Xhold537 data_array.data1\[3\]\[9\] VGND VGND VPWR VPWR net2188 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold548 data_array.data0\[2\]\[0\] VGND VGND VPWR VPWR net2199 sky130_fd_sc_hd__dlygate4sd3_1
X_09950_ net1028 net3622 net377 VGND VGND VPWR VPWR _01699_ sky130_fd_sc_hd__mux2_1
Xhold559 data_array.data0\[13\]\[63\] VGND VGND VPWR VPWR net2210 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08901_ net902 net2678 net437 VGND VGND VPWR VPWR _00658_ sky130_fd_sc_hd__mux2_1
XFILLER_83_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09881_ net945 net4377 net379 VGND VGND VPWR VPWR _01631_ sky130_fd_sc_hd__mux2_1
Xclkbuf_5_12__f_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_5_12__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_170_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08832_ net1895 net916 net447 VGND VGND VPWR VPWR _00590_ sky130_fd_sc_hd__mux2_1
XFILLER_97_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1204 data_array.data1\[3\]\[0\] VGND VGND VPWR VPWR net2855 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1215 data_array.data1\[12\]\[14\] VGND VGND VPWR VPWR net2866 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1226 tag_array.tag0\[12\]\[11\] VGND VGND VPWR VPWR net2877 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1237 data_array.data0\[5\]\[47\] VGND VGND VPWR VPWR net2888 sky130_fd_sc_hd__dlygate4sd3_1
X_05975_ data_array.rdata0\[48\] net1658 net1147 VGND VGND VPWR VPWR _03444_ sky130_fd_sc_hd__o21a_1
Xhold1248 data_array.data1\[11\]\[31\] VGND VGND VPWR VPWR net2899 sky130_fd_sc_hd__dlygate4sd3_1
X_08763_ net771 net3784 net452 VGND VGND VPWR VPWR _00522_ sky130_fd_sc_hd__mux2_1
Xhold1259 data_array.data0\[3\]\[36\] VGND VGND VPWR VPWR net2910 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07714_ net1179 _04925_ _04929_ net1227 VGND VGND VPWR VPWR _04931_ sky130_fd_sc_hd__a22o_1
X_08694_ net2744 net746 net486 VGND VGND VPWR VPWR _00453_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_140_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07645_ data_array.data1\[1\]\[18\] net1534 net1438 data_array.data1\[2\]\[18\] VGND
+ VGND VPWR VPWR _04868_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_101_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07576_ data_array.data1\[0\]\[12\] net1395 net1301 data_array.data1\[3\]\[12\] _04804_
+ VGND VGND VPWR VPWR _04805_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_81_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06527_ _03850_ _03851_ VGND VGND VPWR VPWR _00176_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_24_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09315_ net718 net2356 net546 VGND VGND VPWR VPWR _01069_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_24_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06458_ tag_array.tag0\[4\]\[24\] net1375 net1281 tag_array.tag0\[7\]\[24\] _03788_
+ VGND VGND VPWR VPWR _03789_ sky130_fd_sc_hd__a221o_1
X_09246_ net696 net2369 net647 VGND VGND VPWR VPWR _01000_ sky130_fd_sc_hd__mux2_1
X_09177_ net770 net3880 net629 VGND VGND VPWR VPWR _00931_ sky130_fd_sc_hd__mux2_1
XFILLER_182_839 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06389_ tag_array.tag0\[9\]\[18\] net1565 net1469 tag_array.tag0\[10\]\[18\] VGND
+ VGND VPWR VPWR _03726_ sky130_fd_sc_hd__a22o_1
XFILLER_147_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08128_ data_array.data1\[12\]\[62\] net1415 net1321 data_array.data1\[15\]\[62\]
+ _05306_ VGND VGND VPWR VPWR _05307_ sky130_fd_sc_hd__a221o_1
XFILLER_181_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08059_ data_array.data1\[5\]\[56\] net1533 net1437 data_array.data1\[6\]\[56\] VGND
+ VGND VPWR VPWR _05244_ sky130_fd_sc_hd__a22o_1
X_11070_ net2962 net982 net328 VGND VGND VPWR VPWR _02813_ sky130_fd_sc_hd__mux2_1
XFILLER_0_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_164_3512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_164_3523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput102 mem_rdata[12] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_1
X_10021_ net1000 net2604 net555 VGND VGND VPWR VPWR _01770_ sky130_fd_sc_hd__mux2_1
Xinput113 mem_rdata[22] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_1
XFILLER_89_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput124 mem_rdata[32] VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_1
XFILLER_131_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput135 mem_rdata[42] VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_1
Xhold2450 data_array.data1\[10\]\[7\] VGND VGND VPWR VPWR net4101 sky130_fd_sc_hd__dlygate4sd3_1
Xinput146 mem_rdata[52] VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput157 mem_rdata[62] VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_1
Xhold2461 data_array.data0\[6\]\[44\] VGND VGND VPWR VPWR net4112 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2472 data_array.data0\[3\]\[2\] VGND VGND VPWR VPWR net4123 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2483 data_array.data0\[3\]\[45\] VGND VGND VPWR VPWR net4134 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2494 data_array.data0\[6\]\[33\] VGND VGND VPWR VPWR net4145 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1760 data_array.data0\[6\]\[0\] VGND VGND VPWR VPWR net3411 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1771 data_array.data0\[10\]\[12\] VGND VGND VPWR VPWR net3422 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11972_ clknet_leaf_243_clk _00780_ VGND VGND VPWR VPWR data_array.data0\[4\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1782 data_array.data1\[6\]\[55\] VGND VGND VPWR VPWR net3433 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1793 data_array.data0\[15\]\[6\] VGND VGND VPWR VPWR net3444 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13711_ clknet_leaf_83_clk _02340_ VGND VGND VPWR VPWR data_array.data1\[1\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_647 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10923_ net1049 net2157 net532 VGND VGND VPWR VPWR _02668_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13642_ clknet_leaf_251_clk _02271_ VGND VGND VPWR VPWR data_array.data1\[15\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_10854_ net1071 net2396 net523 VGND VGND VPWR VPWR _02599_ sky130_fd_sc_hd__mux2_1
XFILLER_13_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13573_ clknet_leaf_29_clk _02202_ VGND VGND VPWR VPWR tag_array.dirty1\[1\] sky130_fd_sc_hd__dfxtp_1
X_10785_ net2092 net1090 net505 VGND VGND VPWR VPWR _02530_ sky130_fd_sc_hd__mux2_1
X_12524_ clknet_leaf_195_clk _01218_ VGND VGND VPWR VPWR tag_array.tag1\[11\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12455_ clknet_leaf_81_clk _01149_ VGND VGND VPWR VPWR data_array.data1\[9\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_136_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11406_ clknet_leaf_232_clk _00216_ VGND VGND VPWR VPWR tag_array.tag1\[7\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_125_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12386_ clknet_leaf_71_clk _01080_ VGND VGND VPWR VPWR data_array.data0\[14\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_10_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_1015 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14125_ clknet_leaf_218_clk _02754_ VGND VGND VPWR VPWR data_array.data0\[1\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
X_11337_ net944 net3167 net795 VGND VGND VPWR VPWR _03080_ sky130_fd_sc_hd__mux2_1
XFILLER_126_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14056_ clknet_leaf_265_clk _02685_ VGND VGND VPWR VPWR data_array.data1\[6\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
X_11268_ net958 net3365 net681 VGND VGND VPWR VPWR _03011_ sky130_fd_sc_hd__mux2_1
X_13007_ clknet_leaf_8_clk _01701_ VGND VGND VPWR VPWR data_array.data0\[3\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_37_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10219_ net929 net2827 net355 VGND VGND VPWR VPWR _01966_ sky130_fd_sc_hd__mux2_1
X_11199_ net979 net4362 net656 VGND VGND VPWR VPWR _02942_ sky130_fd_sc_hd__mux2_1
XFILLER_0_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05760_ fsm.tag_out1\[17\] net17 VGND VGND VPWR VPWR _03277_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13909_ clknet_leaf_200_clk _02538_ VGND VGND VPWR VPWR data_array.data1\[4\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05691_ fsm.tag_out0\[7\] net6 VGND VGND VPWR VPWR _03208_ sky130_fd_sc_hd__and2b_1
XFILLER_36_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07430_ data_array.data0\[13\]\[63\] net1556 net1460 data_array.data0\[14\]\[63\]
+ VGND VGND VPWR VPWR _04672_ sky130_fd_sc_hd__a22o_1
XFILLER_50_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07361_ net1192 _04603_ _04607_ net1618 VGND VGND VPWR VPWR _04610_ sky130_fd_sc_hd__a22o_1
X_09100_ net884 net3935 net411 VGND VGND VPWR VPWR _00854_ sky130_fd_sc_hd__mux2_1
X_06312_ tag_array.tag0\[9\]\[11\] net1593 net1497 tag_array.tag0\[10\]\[11\] VGND
+ VGND VPWR VPWR _03656_ sky130_fd_sc_hd__a22o_1
X_07292_ data_array.data0\[12\]\[50\] net1348 net1254 data_array.data0\[15\]\[50\]
+ _04546_ VGND VGND VPWR VPWR _04547_ sky130_fd_sc_hd__a221o_1
X_09031_ net1930 net902 net421 VGND VGND VPWR VPWR _00786_ sky130_fd_sc_hd__mux2_1
X_06243_ tag_array.tag0\[12\]\[5\] net1410 net1316 tag_array.tag0\[15\]\[5\] _03592_
+ VGND VGND VPWR VPWR _03593_ sky130_fd_sc_hd__a221o_1
XFILLER_176_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06174_ net1230 _03521_ net1182 _03529_ VGND VGND VPWR VPWR _03531_ sky130_fd_sc_hd__a22o_1
XFILLER_7_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold301 data_array.data0\[8\]\[11\] VGND VGND VPWR VPWR net1952 sky130_fd_sc_hd__dlygate4sd3_1
Xhold312 data_array.data1\[4\]\[32\] VGND VGND VPWR VPWR net1963 sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 data_array.data1\[1\]\[30\] VGND VGND VPWR VPWR net1974 sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 data_array.data0\[0\]\[5\] VGND VGND VPWR VPWR net1985 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_265_clk clknet_5_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_265_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_105_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold345 data_array.data0\[0\]\[6\] VGND VGND VPWR VPWR net1996 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold356 tag_array.tag1\[4\]\[15\] VGND VGND VPWR VPWR net2007 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold367 data_array.data0\[8\]\[52\] VGND VGND VPWR VPWR net2018 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold378 data_array.data0\[8\]\[41\] VGND VGND VPWR VPWR net2029 sky130_fd_sc_hd__dlygate4sd3_1
Xhold389 data_array.data1\[1\]\[22\] VGND VGND VPWR VPWR net2040 sky130_fd_sc_hd__dlygate4sd3_1
X_09933_ net1096 net4547 net376 VGND VGND VPWR VPWR _01682_ sky130_fd_sc_hd__mux2_1
Xfanout803 net806 VGND VGND VPWR VPWR net803 sky130_fd_sc_hd__buf_2
Xfanout814 net815 VGND VGND VPWR VPWR net814 sky130_fd_sc_hd__buf_2
Xfanout825 _05353_ VGND VGND VPWR VPWR net825 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout847 net853 VGND VGND VPWR VPWR net847 sky130_fd_sc_hd__buf_6
X_09864_ net1012 net4445 net382 VGND VGND VPWR VPWR _01614_ sky130_fd_sc_hd__mux2_1
Xfanout858 net859 VGND VGND VPWR VPWR net858 sky130_fd_sc_hd__clkbuf_2
XFILLER_112_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout869 _05540_ VGND VGND VPWR VPWR net869 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1001 data_array.data1\[15\]\[63\] VGND VGND VPWR VPWR net2652 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1012 data_array.data1\[0\]\[53\] VGND VGND VPWR VPWR net2663 sky130_fd_sc_hd__dlygate4sd3_1
X_08815_ net1856 net986 net446 VGND VGND VPWR VPWR _00573_ sky130_fd_sc_hd__mux2_1
Xhold1023 tag_array.tag1\[15\]\[16\] VGND VGND VPWR VPWR net2674 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_86_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09795_ net1029 net4070 net392 VGND VGND VPWR VPWR _01546_ sky130_fd_sc_hd__mux2_1
Xhold1034 data_array.data0\[2\]\[56\] VGND VGND VPWR VPWR net2685 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1045 data_array.data0\[5\]\[40\] VGND VGND VPWR VPWR net2696 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1056 data_array.data0\[10\]\[30\] VGND VGND VPWR VPWR net2707 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_761 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1067 data_array.data1\[3\]\[2\] VGND VGND VPWR VPWR net2718 sky130_fd_sc_hd__dlygate4sd3_1
X_08746_ net740 net3523 net464 VGND VGND VPWR VPWR _00505_ sky130_fd_sc_hd__mux2_1
X_05958_ data_array.rdata1\[42\] net832 net841 VGND VGND VPWR VPWR _03433_ sky130_fd_sc_hd__a21o_1
Xhold1078 data_array.data1\[8\]\[58\] VGND VGND VPWR VPWR net2729 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1089 tag_array.tag1\[8\]\[9\] VGND VGND VPWR VPWR net2740 sky130_fd_sc_hd__dlygate4sd3_1
X_05889_ data_array.rdata1\[19\] net832 net841 VGND VGND VPWR VPWR _03387_ sky130_fd_sc_hd__a21o_1
X_08677_ net715 net2447 net499 VGND VGND VPWR VPWR _00436_ sky130_fd_sc_hd__mux2_1
XFILLER_26_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07628_ data_array.data1\[13\]\[17\] net1526 net1430 data_array.data1\[14\]\[17\]
+ VGND VGND VPWR VPWR _04852_ sky130_fd_sc_hd__a22o_1
XFILLER_54_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07559_ net1635 _04783_ _04787_ net1209 VGND VGND VPWR VPWR _04790_ sky130_fd_sc_hd__a22o_1
XFILLER_41_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_3382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10570_ net924 net4308 net453 VGND VGND VPWR VPWR _02315_ sky130_fd_sc_hd__mux2_1
XFILLER_139_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_118_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09229_ net762 net2666 net647 VGND VGND VPWR VPWR _00983_ sky130_fd_sc_hd__mux2_1
XFILLER_155_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12240_ clknet_leaf_184_clk _00170_ VGND VGND VPWR VPWR fsm.tag_out1\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_256_clk clknet_5_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_256_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12171_ clknet_leaf_171_clk _00979_ VGND VGND VPWR VPWR tag_array.tag0\[14\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_123_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11122_ net1031 net3739 net551 VGND VGND VPWR VPWR _02865_ sky130_fd_sc_hd__mux2_1
XFILLER_174_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold890 data_array.data1\[7\]\[37\] VGND VGND VPWR VPWR net2541 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11053_ net2143 net1048 net333 VGND VGND VPWR VPWR _02796_ sky130_fd_sc_hd__mux2_1
XFILLER_27_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10004_ net1071 net2987 net564 VGND VGND VPWR VPWR _01753_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2280 data_array.data1\[9\]\[10\] VGND VGND VPWR VPWR net3931 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2291 data_array.data0\[3\]\[60\] VGND VGND VPWR VPWR net3942 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_114_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1590 data_array.data0\[12\]\[2\] VGND VGND VPWR VPWR net3241 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11955_ clknet_leaf_52_clk _00763_ VGND VGND VPWR VPWR data_array.data0\[4\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10906_ net862 net3719 net523 VGND VGND VPWR VPWR _02651_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_177_3758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_177_3769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11886_ clknet_leaf_92_clk _00694_ VGND VGND VPWR VPWR data_array.data0\[5\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_103_Left_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13625_ clknet_leaf_30_clk _02254_ VGND VGND VPWR VPWR data_array.data0\[9\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
X_10837_ net2032 net883 net502 VGND VGND VPWR VPWR _02582_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_82_Right_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13556_ clknet_leaf_5_clk _02185_ VGND VGND VPWR VPWR data_array.data1\[0\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
X_10768_ net900 net4304 net493 VGND VGND VPWR VPWR _02513_ sky130_fd_sc_hd__mux2_1
X_12507_ clknet_leaf_41_clk _01201_ VGND VGND VPWR VPWR data_array.data1\[9\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_173_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13487_ clknet_leaf_181_clk _02117_ VGND VGND VPWR VPWR tag_array.tag0\[15\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_10699_ net2455 net922 net485 VGND VGND VPWR VPWR _02444_ sky130_fd_sc_hd__mux2_1
XFILLER_8_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12438_ clknet_leaf_13_clk _01132_ VGND VGND VPWR VPWR data_array.data0\[14\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_154_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_247_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_247_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_39_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12369_ clknet_leaf_1_clk _00046_ VGND VGND VPWR VPWR data_array.rdata0\[51\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_39_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_112_Left_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14108_ clknet_leaf_126_clk _02737_ VGND VGND VPWR VPWR data_array.data0\[1\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_91_Right_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_566 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14039_ clknet_leaf_64_clk _02668_ VGND VGND VPWR VPWR data_array.data1\[6\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_06930_ data_array.data0\[5\]\[17\] net1528 net1432 data_array.data0\[6\]\[17\] VGND
+ VGND VPWR VPWR _04218_ sky130_fd_sc_hd__a22o_1
XFILLER_80_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06861_ data_array.data0\[0\]\[11\] net1378 net1284 data_array.data0\[3\]\[11\] _04154_
+ VGND VGND VPWR VPWR _04155_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_52_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08600_ net724 net3533 net535 VGND VGND VPWR VPWR _00359_ sky130_fd_sc_hd__mux2_1
X_05812_ _03180_ _03189_ _03205_ _03210_ VGND VGND VPWR VPWR _03329_ sky130_fd_sc_hd__or4_1
X_09580_ net1029 net3572 net400 VGND VGND VPWR VPWR _01332_ sky130_fd_sc_hd__mux2_1
X_06792_ data_array.data0\[9\]\[5\] net1553 net1457 data_array.data0\[10\]\[5\] VGND
+ VGND VPWR VPWR _04092_ sky130_fd_sc_hd__a22o_1
XFILLER_103_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08531_ _05552_ net813 VGND VGND VPWR VPWR _05592_ sky130_fd_sc_hd__nand2b_4
X_05743_ net31 fsm.tag_out1\[1\] VGND VGND VPWR VPWR _03260_ sky130_fd_sc_hd__and2b_1
XFILLER_36_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08462_ net1998 net860 net693 VGND VGND VPWR VPWR _00283_ sky130_fd_sc_hd__mux2_1
X_05674_ _03187_ _03188_ _03189_ _03190_ VGND VGND VPWR VPWR _03191_ sky130_fd_sc_hd__or4_1
X_07413_ data_array.data0\[8\]\[61\] net1361 net1267 data_array.data0\[11\]\[61\]
+ _04656_ VGND VGND VPWR VPWR _04657_ sky130_fd_sc_hd__a221o_1
X_08393_ net2671 net955 net690 VGND VGND VPWR VPWR _00260_ sky130_fd_sc_hd__mux2_1
XFILLER_23_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07344_ data_array.data0\[1\]\[55\] net1534 net1438 data_array.data0\[2\]\[55\] VGND
+ VGND VPWR VPWR _04594_ sky130_fd_sc_hd__a22o_1
XFILLER_177_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07275_ _04530_ _04531_ VGND VGND VPWR VPWR _00042_ sky130_fd_sc_hd__or2_1
XFILLER_128_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09014_ net2141 net971 net418 VGND VGND VPWR VPWR _00769_ sky130_fd_sc_hd__mux2_1
X_06226_ tag_array.tag0\[5\]\[3\] net1561 net1465 tag_array.tag0\[6\]\[3\] VGND VGND
+ VPWR VPWR _03578_ sky130_fd_sc_hd__a22o_1
XFILLER_164_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_152_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_238_clk clknet_5_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_238_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold120 tag_array.tag1\[4\]\[13\] VGND VGND VPWR VPWR net1771 sky130_fd_sc_hd__dlygate4sd3_1
X_06157_ net26 net27 VGND VGND VPWR VPWR _03514_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_76_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold131 data_array.data0\[0\]\[9\] VGND VGND VPWR VPWR net1782 sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 data_array.data0\[4\]\[22\] VGND VGND VPWR VPWR net1793 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold153 data_array.data1\[1\]\[7\] VGND VGND VPWR VPWR net1804 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold164 data_array.data1\[4\]\[29\] VGND VGND VPWR VPWR net1815 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 data_array.data1\[0\]\[44\] VGND VGND VPWR VPWR net1826 sky130_fd_sc_hd__dlygate4sd3_1
X_06088_ data_array.rdata0\[3\] net1140 net1114 data_array.rdata1\[3\] VGND VGND VPWR
+ VPWR net296 sky130_fd_sc_hd__a22o_1
Xhold186 data_array.data0\[8\]\[40\] VGND VGND VPWR VPWR net1837 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout600 net601 VGND VGND VPWR VPWR net600 sky130_fd_sc_hd__buf_4
Xhold197 data_array.data1\[4\]\[14\] VGND VGND VPWR VPWR net1848 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout611 _05576_ VGND VGND VPWR VPWR net611 sky130_fd_sc_hd__buf_4
XFILLER_99_970 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1609 net1612 VGND VGND VPWR VPWR net1609 sky130_fd_sc_hd__clkbuf_4
X_09916_ net744 net3616 net602 VGND VGND VPWR VPWR _01666_ sky130_fd_sc_hd__mux2_1
Xfanout622 _05567_ VGND VGND VPWR VPWR net622 sky130_fd_sc_hd__buf_4
XFILLER_120_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout633 net636 VGND VGND VPWR VPWR net633 sky130_fd_sc_hd__buf_4
Xfanout644 _05557_ VGND VGND VPWR VPWR net644 sky130_fd_sc_hd__clkbuf_4
XFILLER_113_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout655 net660 VGND VGND VPWR VPWR net655 sky130_fd_sc_hd__clkbuf_8
Xfanout666 _05549_ VGND VGND VPWR VPWR net666 sky130_fd_sc_hd__clkbuf_8
Xfanout677 net679 VGND VGND VPWR VPWR net677 sky130_fd_sc_hd__clkbuf_8
XFILLER_101_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09847_ net1080 net3305 net384 VGND VGND VPWR VPWR _01597_ sky130_fd_sc_hd__mux2_1
Xfanout688 net689 VGND VGND VPWR VPWR net688 sky130_fd_sc_hd__buf_4
Xfanout699 _05411_ VGND VGND VPWR VPWR net699 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_160_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09778_ net1097 net2965 net390 VGND VGND VPWR VPWR _01529_ sky130_fd_sc_hd__mux2_1
XFILLER_100_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08729_ net1777 net706 net476 VGND VGND VPWR VPWR _00488_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_159_3411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11740_ clknet_leaf_0_clk _00548_ VGND VGND VPWR VPWR data_array.data0\[8\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11671_ clknet_leaf_167_clk _00479_ VGND VGND VPWR VPWR tag_array.tag1\[1\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_13410_ clknet_leaf_67_clk _02040_ VGND VGND VPWR VPWR data_array.data1\[8\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_169_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10622_ net2253 net974 net467 VGND VGND VPWR VPWR _02367_ sky130_fd_sc_hd__mux2_1
XFILLER_53_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14390_ clknet_leaf_121_clk _03013_ VGND VGND VPWR VPWR data_array.data1\[10\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_12_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13341_ clknet_leaf_25_clk _01971_ VGND VGND VPWR VPWR data_array.data0\[10\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10553_ net995 net3372 net460 VGND VGND VPWR VPWR _02298_ sky130_fd_sc_hd__mux2_1
XFILLER_128_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13272_ clknet_leaf_27_clk _01902_ VGND VGND VPWR VPWR data_array.data0\[11\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
X_10484_ net1009 net2925 net344 VGND VGND VPWR VPWR _02229_ sky130_fd_sc_hd__mux2_1
XFILLER_183_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_229_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_229_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12223_ clknet_leaf_147_clk _00176_ VGND VGND VPWR VPWR fsm.tag_out1\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_907 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12154_ clknet_leaf_164_clk _00962_ VGND VGND VPWR VPWR tag_array.tag0\[13\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_111_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11105_ net1098 net2884 net543 VGND VGND VPWR VPWR _02848_ sky130_fd_sc_hd__mux2_1
XFILLER_151_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12085_ clknet_leaf_36_clk _00893_ VGND VGND VPWR VPWR data_array.data1\[14\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_34_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11036_ net2046 net857 net338 VGND VGND VPWR VPWR _02780_ sky130_fd_sc_hd__mux2_1
XFILLER_110_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_804 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12987_ clknet_leaf_247_clk _01681_ VGND VGND VPWR VPWR data_array.data0\[3\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_73_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11938_ clknet_leaf_94_clk _00746_ VGND VGND VPWR VPWR data_array.data0\[4\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_222 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11869_ clknet_leaf_104_clk _00677_ VGND VGND VPWR VPWR data_array.data0\[5\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13608_ clknet_leaf_89_clk _02237_ VGND VGND VPWR VPWR data_array.data0\[9\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_159_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13539_ clknet_leaf_117_clk _02168_ VGND VGND VPWR VPWR data_array.data1\[0\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_31_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07060_ data_array.data0\[9\]\[29\] net1570 net1474 data_array.data0\[10\]\[29\]
+ VGND VGND VPWR VPWR _04336_ sky130_fd_sc_hd__a22o_1
XFILLER_134_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_120_Left_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06011_ data_array.rdata0\[60\] net1659 net1149 VGND VGND VPWR VPWR _03468_ sky130_fd_sc_hd__o21a_1
XFILLER_161_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput203 net203 VGND VGND VPWR VPWR cpu_rdata[44] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_93_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput214 net214 VGND VGND VPWR VPWR cpu_rdata[54] sky130_fd_sc_hd__clkbuf_4
XFILLER_114_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput225 net225 VGND VGND VPWR VPWR cpu_rdata[6] sky130_fd_sc_hd__buf_4
Xoutput236 net236 VGND VGND VPWR VPWR mem_addr[15] sky130_fd_sc_hd__buf_2
Xoutput247 net247 VGND VGND VPWR VPWR mem_addr[25] sky130_fd_sc_hd__buf_2
XFILLER_114_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput258 net258 VGND VGND VPWR VPWR mem_addr[6] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput269 net269 VGND VGND VPWR VPWR mem_wdata[15] sky130_fd_sc_hd__buf_2
X_07962_ data_array.data1\[13\]\[47\] net1588 net1492 data_array.data1\[14\]\[47\]
+ VGND VGND VPWR VPWR _05156_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_71_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09701_ net784 net3420 net609 VGND VGND VPWR VPWR _01453_ sky130_fd_sc_hd__mux2_1
X_06913_ data_array.data0\[9\]\[16\] net1548 net1452 data_array.data0\[10\]\[16\]
+ VGND VGND VPWR VPWR _04202_ sky130_fd_sc_hd__a22o_1
X_07893_ data_array.data1\[8\]\[41\] net1335 net1241 data_array.data1\[11\]\[41\]
+ _05092_ VGND VGND VPWR VPWR _05093_ sky130_fd_sc_hd__a221o_1
XFILLER_67_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09632_ net761 net4435 net617 VGND VGND VPWR VPWR _01384_ sky130_fd_sc_hd__mux2_1
X_06844_ net1630 _04133_ _04137_ net1204 VGND VGND VPWR VPWR _04140_ sky130_fd_sc_hd__a22o_1
XFILLER_167_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09563_ net1097 net4457 net398 VGND VGND VPWR VPWR _01315_ sky130_fd_sc_hd__mux2_1
X_06775_ data_array.data0\[8\]\[3\] net1377 net1283 data_array.data0\[11\]\[3\] _04076_
+ VGND VGND VPWR VPWR _04077_ sky130_fd_sc_hd__a221o_1
XFILLER_24_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08514_ _03514_ _03527_ VGND VGND VPWR VPWR _05580_ sky130_fd_sc_hd__nor2_1
XFILLER_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05726_ net18 fsm.tag_out1\[18\] VGND VGND VPWR VPWR _03243_ sky130_fd_sc_hd__nand2b_1
X_09494_ net753 net4000 net625 VGND VGND VPWR VPWR _01247_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_137_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08445_ net151 net86 net1643 VGND VGND VPWR VPWR _05533_ sky130_fd_sc_hd__mux2_1
X_05657_ net4 fsm.tag_out0\[5\] VGND VGND VPWR VPWR _03174_ sky130_fd_sc_hd__and2b_1
XFILLER_23_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_154_3330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08376_ net126 net61 net1638 VGND VGND VPWR VPWR _05487_ sky130_fd_sc_hd__mux2_1
X_07327_ data_array.data0\[4\]\[53\] net1332 net1238 data_array.data0\[7\]\[53\] _04578_
+ VGND VGND VPWR VPWR _04579_ sky130_fd_sc_hd__a221o_1
XFILLER_20_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_150_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07258_ data_array.data0\[13\]\[47\] net1577 net1481 data_array.data0\[14\]\[47\]
+ VGND VGND VPWR VPWR _04516_ sky130_fd_sc_hd__a22o_1
XFILLER_180_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06209_ tag_array.tag0\[9\]\[2\] net1559 net1464 tag_array.tag0\[10\]\[2\] VGND VGND
+ VPWR VPWR _03562_ sky130_fd_sc_hd__a22o_1
X_07189_ data_array.data0\[8\]\[41\] net1337 net1243 data_array.data0\[11\]\[41\]
+ _04452_ VGND VGND VPWR VPWR _04453_ sky130_fd_sc_hd__a221o_1
XFILLER_133_820 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1406 net1422 VGND VGND VPWR VPWR net1406 sky130_fd_sc_hd__buf_2
Xfanout1417 net1421 VGND VGND VPWR VPWR net1417 sky130_fd_sc_hd__clkbuf_4
Xfanout1428 net1447 VGND VGND VPWR VPWR net1428 sky130_fd_sc_hd__buf_2
Xfanout430 net431 VGND VGND VPWR VPWR net430 sky130_fd_sc_hd__buf_4
Xfanout441 _05608_ VGND VGND VPWR VPWR net441 sky130_fd_sc_hd__clkbuf_8
Xfanout1439 net1440 VGND VGND VPWR VPWR net1439 sky130_fd_sc_hd__clkbuf_4
XFILLER_24_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout452 _05606_ VGND VGND VPWR VPWR net452 sky130_fd_sc_hd__buf_2
Xfanout463 net464 VGND VGND VPWR VPWR net463 sky130_fd_sc_hd__buf_4
XFILLER_87_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout474 net477 VGND VGND VPWR VPWR net474 sky130_fd_sc_hd__clkbuf_4
Xfanout485 net486 VGND VGND VPWR VPWR net485 sky130_fd_sc_hd__clkbuf_4
XFILLER_24_1057 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout496 net499 VGND VGND VPWR VPWR net496 sky130_fd_sc_hd__clkbuf_8
XFILLER_111_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12910_ clknet_leaf_51_clk _01604_ VGND VGND VPWR VPWR data_array.data0\[13\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_100_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13890_ clknet_leaf_202_clk _02519_ VGND VGND VPWR VPWR data_array.data1\[3\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_859 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12841_ clknet_leaf_60_clk _01535_ VGND VGND VPWR VPWR data_array.data0\[12\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_126_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12772_ clknet_leaf_165_clk _01466_ VGND VGND VPWR VPWR tag_array.tag0\[6\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_174_3706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ clknet_leaf_173_clk _00531_ VGND VGND VPWR VPWR tag_array.tag0\[9\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14442_ clknet_leaf_254_clk _03065_ VGND VGND VPWR VPWR data_array.data1\[7\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11654_ clknet_leaf_234_clk _00462_ VGND VGND VPWR VPWR tag_array.tag1\[2\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_10605_ net1833 net1040 net466 VGND VGND VPWR VPWR _02350_ sky130_fd_sc_hd__mux2_1
X_14373_ clknet_leaf_204_clk _02996_ VGND VGND VPWR VPWR data_array.data1\[10\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_11585_ clknet_leaf_167_clk _00393_ VGND VGND VPWR VPWR tag_array.tag1\[4\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_80_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13324_ clknet_leaf_89_clk _01954_ VGND VGND VPWR VPWR data_array.data0\[10\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10536_ net1062 net4294 net462 VGND VGND VPWR VPWR _02281_ sky130_fd_sc_hd__mux2_1
XFILLER_156_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13255_ clknet_leaf_31_clk _01885_ VGND VGND VPWR VPWR data_array.data0\[11\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_108_Right_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10467_ net1077 net2682 net345 VGND VGND VPWR VPWR _02212_ sky130_fd_sc_hd__mux2_1
X_12206_ clknet_leaf_147_clk _00135_ VGND VGND VPWR VPWR fsm.tag_out0\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_159_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13186_ clknet_leaf_201_clk _00079_ VGND VGND VPWR VPWR data_array.rdata1\[23\] sky130_fd_sc_hd__dfxtp_1
X_10398_ net1989 net1062 net669 VGND VGND VPWR VPWR _02144_ sky130_fd_sc_hd__mux2_1
XFILLER_69_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12137_ clknet_leaf_160_clk _00945_ VGND VGND VPWR VPWR tag_array.tag0\[12\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_12068_ clknet_leaf_42_clk _00876_ VGND VGND VPWR VPWR data_array.data1\[14\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_65_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11019_ net1924 net926 net336 VGND VGND VPWR VPWR _02763_ sky130_fd_sc_hd__mux2_1
XFILLER_38_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06560_ _03880_ _03881_ VGND VGND VPWR VPWR _00179_ sky130_fd_sc_hd__or2_1
X_06491_ tag_array.tag1\[0\]\[2\] net1351 net1257 tag_array.tag1\[3\]\[2\] _03818_
+ VGND VGND VPWR VPWR _03819_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_47_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08230_ net1651 net1158 net11 VGND VGND VPWR VPWR _05388_ sky130_fd_sc_hd__and3_1
XFILLER_166_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08161_ tag_array.dirty0\[8\] net1403 net1309 tag_array.dirty0\[11\] _05336_ VGND
+ VGND VPWR VPWR _05337_ sky130_fd_sc_hd__a221o_1
X_07112_ data_array.data0\[12\]\[34\] net1340 net1246 data_array.data0\[15\]\[34\]
+ _04382_ VGND VGND VPWR VPWR _04383_ sky130_fd_sc_hd__a221o_1
XFILLER_118_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08092_ data_array.data1\[1\]\[59\] net1572 net1476 data_array.data1\[2\]\[59\] VGND
+ VGND VPWR VPWR _05274_ sky130_fd_sc_hd__a22o_1
XFILLER_173_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07043_ net1222 _04315_ _04319_ net1173 VGND VGND VPWR VPWR _04321_ sky130_fd_sc_hd__a22o_1
Xclkload40 clknet_leaf_20_clk VGND VGND VPWR VPWR clkload40/X sky130_fd_sc_hd__clkbuf_4
XFILLER_146_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload51 clknet_leaf_249_clk VGND VGND VPWR VPWR clkload51/X sky130_fd_sc_hd__clkbuf_4
Xclkload62 clknet_leaf_29_clk VGND VGND VPWR VPWR clkload62/Y sky130_fd_sc_hd__inv_6
Xclkload73 clknet_leaf_239_clk VGND VGND VPWR VPWR clkload73/Y sky130_fd_sc_hd__inv_12
XFILLER_161_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload84 clknet_leaf_44_clk VGND VGND VPWR VPWR clkload84/Y sky130_fd_sc_hd__clkinv_8
Xclkload95 clknet_leaf_57_clk VGND VGND VPWR VPWR clkload95/Y sky130_fd_sc_hd__bufinv_16
XFILLER_102_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2802 data_array.data0\[3\]\[18\] VGND VGND VPWR VPWR net4453 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_141_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08994_ net1737 net1048 net422 VGND VGND VPWR VPWR _00749_ sky130_fd_sc_hd__mux2_1
Xhold2813 data_array.data1\[2\]\[43\] VGND VGND VPWR VPWR net4464 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2824 data_array.data1\[14\]\[33\] VGND VGND VPWR VPWR net4475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2835 data_array.data1\[6\]\[59\] VGND VGND VPWR VPWR net4486 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2846 data_array.data0\[11\]\[44\] VGND VGND VPWR VPWR net4497 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07945_ net1217 _05135_ _05139_ net1169 VGND VGND VPWR VPWR _05141_ sky130_fd_sc_hd__a22o_1
Xhold2857 data_array.data0\[11\]\[30\] VGND VGND VPWR VPWR net4508 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2868 data_array.data1\[11\]\[48\] VGND VGND VPWR VPWR net4519 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2879 data_array.data1\[6\]\[23\] VGND VGND VPWR VPWR net4530 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07876_ data_array.data1\[5\]\[39\] net1539 net1443 data_array.data1\[6\]\[39\] VGND
+ VGND VPWR VPWR _05078_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_3_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09615_ net888 net3885 net395 VGND VGND VPWR VPWR _01367_ sky130_fd_sc_hd__mux2_1
X_06827_ data_array.data0\[5\]\[8\] net1534 net1438 data_array.data0\[6\]\[8\] VGND
+ VGND VPWR VPWR _04124_ sky130_fd_sc_hd__a22o_1
XFILLER_84_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09546_ net745 net3678 net618 VGND VGND VPWR VPWR _01299_ sky130_fd_sc_hd__mux2_1
X_06758_ _04060_ _04061_ VGND VGND VPWR VPWR _00011_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_104_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05709_ _03219_ _03222_ _03223_ _03225_ VGND VGND VPWR VPWR _03226_ sky130_fd_sc_hd__or4_1
X_09477_ net718 net3285 net654 VGND VGND VPWR VPWR _01230_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_84_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06689_ tag_array.tag1\[4\]\[20\] net1349 net1255 tag_array.tag1\[7\]\[20\] _03998_
+ VGND VGND VPWR VPWR _03999_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_84_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_121_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08428_ net1123 _05521_ VGND VGND VPWR VPWR _05522_ sky130_fd_sc_hd__and2_1
XFILLER_140_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload1 clknet_5_3__leaf_clk VGND VGND VPWR VPWR clkload1/X sky130_fd_sc_hd__clkbuf_8
XFILLER_184_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08359_ net1124 _05475_ VGND VGND VPWR VPWR _05476_ sky130_fd_sc_hd__and2_1
X_11370_ net1646 net4261 net619 VGND VGND VPWR VPWR _03113_ sky130_fd_sc_hd__mux2_1
XFILLER_138_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10321_ net2729 net878 net637 VGND VGND VPWR VPWR _02068_ sky130_fd_sc_hd__mux2_1
XFILLER_30_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13040_ clknet_leaf_13_clk _01734_ VGND VGND VPWR VPWR data_array.data0\[3\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_124_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10252_ net735 net3790 net595 VGND VGND VPWR VPWR _01999_ sky130_fd_sc_hd__mux2_1
XFILLER_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_167_3565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_3576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10183_ net1073 net3050 net358 VGND VGND VPWR VPWR _01930_ sky130_fd_sc_hd__mux2_1
Xfanout1203 net1212 VGND VGND VPWR VPWR net1203 sky130_fd_sc_hd__buf_4
Xfanout1214 net1215 VGND VGND VPWR VPWR net1214 sky130_fd_sc_hd__buf_4
XFILLER_78_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1225 net1234 VGND VGND VPWR VPWR net1225 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_184_3890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1236 net1237 VGND VGND VPWR VPWR net1236 sky130_fd_sc_hd__clkbuf_4
XFILLER_94_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1247 net1248 VGND VGND VPWR VPWR net1247 sky130_fd_sc_hd__clkbuf_4
XFILLER_78_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1258 net1282 VGND VGND VPWR VPWR net1258 sky130_fd_sc_hd__buf_2
Xfanout1269 net1270 VGND VGND VPWR VPWR net1269 sky130_fd_sc_hd__clkbuf_2
XFILLER_8_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13942_ clknet_leaf_261_clk _02571_ VGND VGND VPWR VPWR data_array.data1\[4\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13873_ clknet_leaf_257_clk _02502_ VGND VGND VPWR VPWR data_array.data1\[3\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12824_ clknet_leaf_129_clk _01518_ VGND VGND VPWR VPWR tag_array.tag1\[0\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12755_ clknet_leaf_108_clk _01449_ VGND VGND VPWR VPWR tag_array.tag0\[5\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_586 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11706_ clknet_leaf_196_clk _00514_ VGND VGND VPWR VPWR tag_array.tag1\[15\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_12686_ clknet_leaf_178_clk _01380_ VGND VGND VPWR VPWR tag_array.tag0\[8\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_14425_ clknet_leaf_57_clk _03048_ VGND VGND VPWR VPWR data_array.data1\[7\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_11637_ clknet_leaf_192_clk _00445_ VGND VGND VPWR VPWR tag_array.tag1\[2\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_156_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14356_ clknet_leaf_268_clk _02979_ VGND VGND VPWR VPWR data_array.data1\[10\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_42_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11568_ clknet_leaf_127_clk _00376_ VGND VGND VPWR VPWR tag_array.tag1\[5\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold708 tag_array.tag1\[8\]\[4\] VGND VGND VPWR VPWR net2359 sky130_fd_sc_hd__dlygate4sd3_1
X_13307_ clknet_leaf_224_clk _01937_ VGND VGND VPWR VPWR data_array.data0\[10\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_116_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10519_ net869 net2535 net351 VGND VGND VPWR VPWR _02264_ sky130_fd_sc_hd__mux2_1
XFILLER_155_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold719 tag_array.tag1\[0\]\[12\] VGND VGND VPWR VPWR net2370 sky130_fd_sc_hd__dlygate4sd3_1
X_14287_ clknet_leaf_81_clk _02916_ VGND VGND VPWR VPWR data_array.data1\[11\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_90_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11499_ clknet_leaf_172_clk _00307_ VGND VGND VPWR VPWR tag_array.valid1\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_90_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13238_ clknet_leaf_45_clk _01868_ VGND VGND VPWR VPWR data_array.data0\[11\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_170_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13169_ clknet_leaf_269_clk _00124_ VGND VGND VPWR VPWR data_array.rdata1\[6\] sky130_fd_sc_hd__dfxtp_1
Xhold2109 data_array.data1\[9\]\[15\] VGND VGND VPWR VPWR net3760 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_3_991 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05991_ data_array.rdata1\[53\] net828 net837 VGND VGND VPWR VPWR _03455_ sky130_fd_sc_hd__a21o_1
Xhold1408 data_array.data0\[5\]\[55\] VGND VGND VPWR VPWR net3059 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1419 data_array.data1\[4\]\[61\] VGND VGND VPWR VPWR net3070 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07730_ data_array.data1\[4\]\[26\] net1335 net1241 data_array.data1\[7\]\[26\] _04944_
+ VGND VGND VPWR VPWR _04945_ sky130_fd_sc_hd__a221o_1
XFILLER_84_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_88_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_751 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07661_ data_array.data1\[13\]\[20\] net1610 net1514 data_array.data1\[14\]\[20\]
+ VGND VGND VPWR VPWR _04882_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_49_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09400_ net1066 net3220 net590 VGND VGND VPWR VPWR _01153_ sky130_fd_sc_hd__mux2_1
X_06612_ tag_array.tag1\[0\]\[13\] net1421 net1327 tag_array.tag1\[3\]\[13\] _03928_
+ VGND VGND VPWR VPWR _03929_ sky130_fd_sc_hd__a221o_1
XFILLER_25_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07592_ net1196 _04813_ _04817_ net1622 VGND VGND VPWR VPWR _04820_ sky130_fd_sc_hd__a22o_1
XFILLER_34_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09331_ net1077 net3454 net403 VGND VGND VPWR VPWR _01084_ sky130_fd_sc_hd__mux2_1
X_06543_ tag_array.tag1\[13\]\[7\] net1611 net1515 tag_array.tag1\[14\]\[7\] VGND
+ VGND VPWR VPWR _03866_ sky130_fd_sc_hd__a22o_1
XFILLER_34_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09262_ net731 net3460 net575 VGND VGND VPWR VPWR _01016_ sky130_fd_sc_hd__mux2_1
X_06474_ tag_array.tag1\[12\]\[1\] net1370 net1276 tag_array.tag1\[15\]\[1\] _03802_
+ VGND VGND VPWR VPWR _03803_ sky130_fd_sc_hd__a221o_1
X_08213_ fsm.tag_out1\[6\] net816 net808 fsm.tag_out0\[6\] _05376_ VGND VGND VPWR
+ VPWR _05377_ sky130_fd_sc_hd__a221o_2
XFILLER_53_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09193_ net708 net3830 net628 VGND VGND VPWR VPWR _00947_ sky130_fd_sc_hd__mux2_1
X_08144_ _05320_ _05321_ VGND VGND VPWR VPWR _00123_ sky130_fd_sc_hd__or2_1
XFILLER_101_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload140 clknet_leaf_222_clk VGND VGND VPWR VPWR clkload140/Y sky130_fd_sc_hd__inv_6
XFILLER_174_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08075_ data_array.data1\[4\]\[57\] net1338 net1244 data_array.data1\[7\]\[57\] _05258_
+ VGND VGND VPWR VPWR _05259_ sky130_fd_sc_hd__a221o_1
Xclkload151 clknet_leaf_228_clk VGND VGND VPWR VPWR clkload151/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload162 clknet_leaf_175_clk VGND VGND VPWR VPWR clkload162/Y sky130_fd_sc_hd__clkinv_2
Xclkload173 clknet_leaf_198_clk VGND VGND VPWR VPWR clkload173/Y sky130_fd_sc_hd__inv_6
X_07026_ data_array.data0\[4\]\[26\] net1338 net1244 data_array.data0\[7\]\[26\] _04304_
+ VGND VGND VPWR VPWR _04305_ sky130_fd_sc_hd__a221o_1
Xclkload184 clknet_leaf_185_clk VGND VGND VPWR VPWR clkload184/Y sky130_fd_sc_hd__clkinv_2
Xclkload195 clknet_leaf_104_clk VGND VGND VPWR VPWR clkload195/Y sky130_fd_sc_hd__clkinv_4
XFILLER_1_939 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2610 tag_array.dirty0\[0\] VGND VGND VPWR VPWR net4261 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2621 tag_array.tag1\[11\]\[21\] VGND VGND VPWR VPWR net4272 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2632 data_array.data0\[3\]\[41\] VGND VGND VPWR VPWR net4283 sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ net856 net3926 net429 VGND VGND VPWR VPWR _00733_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_145_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2643 data_array.data1\[15\]\[12\] VGND VGND VPWR VPWR net4294 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_145_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold46 tag_array.valid1\[12\] VGND VGND VPWR VPWR net1697 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2654 data_array.data0\[7\]\[14\] VGND VGND VPWR VPWR net4305 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1920 data_array.data1\[6\]\[33\] VGND VGND VPWR VPWR net3571 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2665 tag_array.tag1\[5\]\[14\] VGND VGND VPWR VPWR net4316 sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ data_array.data1\[0\]\[44\] net1398 net1304 data_array.data1\[3\]\[44\] _05124_
+ VGND VGND VPWR VPWR _05125_ sky130_fd_sc_hd__a221o_1
Xhold57 tag_array.valid1\[7\] VGND VGND VPWR VPWR net1708 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1931 data_array.data1\[5\]\[29\] VGND VGND VPWR VPWR net3582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2676 tag_array.tag0\[0\]\[23\] VGND VGND VPWR VPWR net4327 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1942 data_array.data0\[12\]\[56\] VGND VGND VPWR VPWR net3593 sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 tag_array.valid0\[1\] VGND VGND VPWR VPWR net1719 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2687 data_array.data1\[6\]\[18\] VGND VGND VPWR VPWR net4338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 data_array.data1\[1\]\[9\] VGND VGND VPWR VPWR net1730 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1953 data_array.data1\[6\]\[30\] VGND VGND VPWR VPWR net3604 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_162_3484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2698 data_array.data1\[12\]\[59\] VGND VGND VPWR VPWR net4349 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1964 data_array.data0\[9\]\[43\] VGND VGND VPWR VPWR net3615 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1975 data_array.data0\[13\]\[16\] VGND VGND VPWR VPWR net3626 sky130_fd_sc_hd__dlygate4sd3_1
X_07859_ data_array.data1\[9\]\[38\] net1588 net1492 data_array.data1\[10\]\[38\]
+ VGND VGND VPWR VPWR _05062_ sky130_fd_sc_hd__a22o_1
XFILLER_45_12 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1986 tag_array.tag0\[8\]\[24\] VGND VGND VPWR VPWR net3637 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1997 tag_array.tag1\[13\]\[10\] VGND VGND VPWR VPWR net3648 sky130_fd_sc_hd__dlygate4sd3_1
X_10870_ net1004 net3494 net515 VGND VGND VPWR VPWR _02615_ sky130_fd_sc_hd__mux2_1
XFILLER_43_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09529_ net712 net2358 net621 VGND VGND VPWR VPWR _01282_ sky130_fd_sc_hd__mux2_1
X_12540_ clknet_leaf_196_clk _01234_ VGND VGND VPWR VPWR tag_array.tag1\[11\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_61_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_84 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12471_ clknet_leaf_194_clk _01165_ VGND VGND VPWR VPWR data_array.data1\[9\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_61_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14210_ clknet_leaf_208_clk _02839_ VGND VGND VPWR VPWR data_array.data0\[2\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
X_11422_ clknet_leaf_45_clk _00232_ VGND VGND VPWR VPWR data_array.data0\[0\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_169_3605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14141_ clknet_leaf_2_clk _02770_ VGND VGND VPWR VPWR data_array.data0\[1\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_169_3616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11353_ net883 net3820 net795 VGND VGND VPWR VPWR _03096_ sky130_fd_sc_hd__mux2_1
X_10304_ net2062 net944 net633 VGND VGND VPWR VPWR _02051_ sky130_fd_sc_hd__mux2_1
X_14072_ clknet_leaf_71_clk _02701_ VGND VGND VPWR VPWR data_array.data1\[6\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11284_ net892 net3699 net674 VGND VGND VPWR VPWR _03027_ sky130_fd_sc_hd__mux2_1
XFILLER_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13023_ clknet_leaf_88_clk _01717_ VGND VGND VPWR VPWR data_array.data0\[3\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
X_10235_ net867 net3502 net356 VGND VGND VPWR VPWR _01982_ sky130_fd_sc_hd__mux2_1
Xfanout1000 _05474_ VGND VGND VPWR VPWR net1000 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_182_3849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1011 _05470_ VGND VGND VPWR VPWR net1011 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1022 net1023 VGND VGND VPWR VPWR net1022 sky130_fd_sc_hd__clkbuf_2
Xfanout1033 _05458_ VGND VGND VPWR VPWR net1033 sky130_fd_sc_hd__dlymetal6s2s_1
X_10166_ net880 net4233 net365 VGND VGND VPWR VPWR _01914_ sky130_fd_sc_hd__mux2_1
Xfanout1044 _05452_ VGND VGND VPWR VPWR net1044 sky130_fd_sc_hd__clkbuf_2
Xfanout1055 _05448_ VGND VGND VPWR VPWR net1055 sky130_fd_sc_hd__buf_1
Xfanout1066 net1067 VGND VGND VPWR VPWR net1066 sky130_fd_sc_hd__clkbuf_2
Xfanout1077 _05436_ VGND VGND VPWR VPWR net1077 sky130_fd_sc_hd__buf_1
XFILLER_120_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1088 net1089 VGND VGND VPWR VPWR net1088 sky130_fd_sc_hd__clkbuf_2
X_10097_ net2749 net737 net638 VGND VGND VPWR VPWR _01846_ sky130_fd_sc_hd__mux2_1
XFILLER_19_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1099 _05426_ VGND VGND VPWR VPWR net1099 sky130_fd_sc_hd__dlymetal6s2s_1
X_13925_ clknet_leaf_40_clk _02554_ VGND VGND VPWR VPWR data_array.data1\[4\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_142_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13856_ clknet_leaf_91_clk _02485_ VGND VGND VPWR VPWR data_array.data1\[3\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12807_ clknet_leaf_98_clk _01501_ VGND VGND VPWR VPWR tag_array.tag1\[0\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_13787_ clknet_leaf_66_clk _02416_ VGND VGND VPWR VPWR data_array.data1\[2\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_10999_ net2082 net1007 net339 VGND VGND VPWR VPWR _02743_ sky130_fd_sc_hd__mux2_1
XFILLER_43_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12738_ clknet_leaf_179_clk _01432_ VGND VGND VPWR VPWR tag_array.tag0\[5\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_26_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12669_ clknet_leaf_4_clk _01363_ VGND VGND VPWR VPWR data_array.data0\[15\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_61_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14408_ clknet_leaf_202_clk _03031_ VGND VGND VPWR VPWR data_array.data1\[10\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
X_06190_ tag_array.tag0\[4\]\[0\] net1405 net1311 tag_array.tag0\[7\]\[0\] _03544_
+ VGND VGND VPWR VPWR _03545_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_160_Right_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14339_ clknet_leaf_41_clk _02968_ VGND VGND VPWR VPWR data_array.data1\[11\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold505 tag_array.tag1\[2\]\[4\] VGND VGND VPWR VPWR net2156 sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 data_array.data0\[4\]\[59\] VGND VGND VPWR VPWR net2167 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold527 data_array.data0\[4\]\[3\] VGND VGND VPWR VPWR net2178 sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 data_array.data1\[12\]\[17\] VGND VGND VPWR VPWR net2189 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold549 data_array.data0\[4\]\[43\] VGND VGND VPWR VPWR net2200 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08900_ net904 net4394 net434 VGND VGND VPWR VPWR _00657_ sky130_fd_sc_hd__mux2_1
X_09880_ net948 net3532 net384 VGND VGND VPWR VPWR _01630_ sky130_fd_sc_hd__mux2_1
XFILLER_170_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08831_ net2118 net920 net446 VGND VGND VPWR VPWR _00589_ sky130_fd_sc_hd__mux2_1
XFILLER_170_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1205 tag_array.tag0\[2\]\[1\] VGND VGND VPWR VPWR net2856 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1216 tag_array.tag1\[12\]\[6\] VGND VGND VPWR VPWR net2867 sky130_fd_sc_hd__dlygate4sd3_1
X_08762_ net777 net3861 net450 VGND VGND VPWR VPWR _00521_ sky130_fd_sc_hd__mux2_1
Xhold1227 tag_array.tag0\[10\]\[0\] VGND VGND VPWR VPWR net2878 sky130_fd_sc_hd__dlygate4sd3_1
X_05974_ net140 net1156 _03442_ _03443_ VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__a22o_1
Xhold1238 data_array.data1\[10\]\[27\] VGND VGND VPWR VPWR net2889 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1249 data_array.data0\[11\]\[2\] VGND VGND VPWR VPWR net2900 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07713_ net1205 _04923_ _04927_ net1631 VGND VGND VPWR VPWR _04930_ sky130_fd_sc_hd__a22o_1
XFILLER_66_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08693_ net2182 net750 net488 VGND VGND VPWR VPWR _00452_ sky130_fd_sc_hd__mux2_1
XFILLER_81_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07644_ data_array.data1\[12\]\[18\] net1383 net1289 data_array.data1\[15\]\[18\]
+ _04866_ VGND VGND VPWR VPWR _04867_ sky130_fd_sc_hd__a221o_1
XFILLER_25_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07575_ data_array.data1\[1\]\[12\] net1586 net1490 data_array.data1\[2\]\[12\] VGND
+ VGND VPWR VPWR _04804_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_81_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09314_ net725 net3023 net551 VGND VGND VPWR VPWR _01068_ sky130_fd_sc_hd__mux2_1
X_06526_ net1232 _03845_ _03849_ net1184 VGND VGND VPWR VPWR _03851_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_24_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09245_ net698 net2610 net646 VGND VGND VPWR VPWR _00999_ sky130_fd_sc_hd__mux2_1
X_06457_ tag_array.tag0\[5\]\[24\] net1562 net1466 tag_array.tag0\[6\]\[24\] VGND
+ VGND VPWR VPWR _03788_ sky130_fd_sc_hd__a22o_1
X_09176_ net776 net4022 net627 VGND VGND VPWR VPWR _00930_ sky130_fd_sc_hd__mux2_1
X_06388_ tag_array.tag0\[0\]\[18\] net1374 net1280 tag_array.tag0\[3\]\[18\] _03724_
+ VGND VGND VPWR VPWR _03725_ sky130_fd_sc_hd__a221o_1
XFILLER_108_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08127_ data_array.data1\[13\]\[62\] net1605 net1509 data_array.data1\[14\]\[62\]
+ VGND VGND VPWR VPWR _05306_ sky130_fd_sc_hd__a22o_1
XFILLER_108_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08058_ data_array.data1\[12\]\[56\] net1341 net1247 data_array.data1\[15\]\[56\]
+ _05242_ VGND VGND VPWR VPWR _05243_ sky130_fd_sc_hd__a221o_1
XFILLER_116_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07009_ net1203 _04283_ _04287_ net1629 VGND VGND VPWR VPWR _04290_ sky130_fd_sc_hd__a22o_1
XFILLER_0_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_164_3513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_24 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_758 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10020_ net1004 net3043 net555 VGND VGND VPWR VPWR _01769_ sky130_fd_sc_hd__mux2_1
XFILLER_103_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput103 mem_rdata[13] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_1
Xinput114 mem_rdata[23] VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__buf_1
XFILLER_102_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput125 mem_rdata[33] VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2440 data_array.data0\[6\]\[1\] VGND VGND VPWR VPWR net4091 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput136 mem_rdata[43] VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_1
XFILLER_130_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2451 data_array.data1\[10\]\[44\] VGND VGND VPWR VPWR net4102 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput147 mem_rdata[53] VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_1
Xinput158 mem_rdata[63] VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2462 data_array.data0\[7\]\[42\] VGND VGND VPWR VPWR net4113 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2473 data_array.data1\[11\]\[4\] VGND VGND VPWR VPWR net4124 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2484 data_array.data1\[15\]\[48\] VGND VGND VPWR VPWR net4135 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1750 data_array.data1\[15\]\[15\] VGND VGND VPWR VPWR net3401 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2495 data_array.data0\[9\]\[39\] VGND VGND VPWR VPWR net4146 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1761 tag_array.tag1\[15\]\[17\] VGND VGND VPWR VPWR net3412 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_5_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11971_ clknet_leaf_20_clk _00779_ VGND VGND VPWR VPWR data_array.data0\[4\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1772 tag_array.tag1\[9\]\[4\] VGND VGND VPWR VPWR net3423 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_99_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1783 data_array.data0\[9\]\[54\] VGND VGND VPWR VPWR net3434 sky130_fd_sc_hd__dlygate4sd3_1
X_13710_ clknet_leaf_268_clk _02339_ VGND VGND VPWR VPWR data_array.data1\[1\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1794 tag_array.tag0\[14\]\[22\] VGND VGND VPWR VPWR net3445 sky130_fd_sc_hd__dlygate4sd3_1
X_10922_ net1054 net4557 net531 VGND VGND VPWR VPWR _02667_ sky130_fd_sc_hd__mux2_1
XFILLER_17_659 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13641_ clknet_leaf_264_clk _02270_ VGND VGND VPWR VPWR data_array.data1\[15\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_10853_ net1074 net3895 net520 VGND VGND VPWR VPWR _02598_ sky130_fd_sc_hd__mux2_1
XFILLER_25_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13572_ clknet_leaf_29_clk _02201_ VGND VGND VPWR VPWR tag_array.dirty1\[2\] sky130_fd_sc_hd__dfxtp_1
X_10784_ net1902 net1094 net508 VGND VGND VPWR VPWR _02529_ sky130_fd_sc_hd__mux2_1
XFILLER_24_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12523_ clknet_leaf_135_clk _01217_ VGND VGND VPWR VPWR tag_array.tag1\[11\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_158_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12454_ clknet_leaf_268_clk _01148_ VGND VGND VPWR VPWR data_array.data1\[9\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11405_ clknet_leaf_98_clk _00215_ VGND VGND VPWR VPWR tag_array.tag1\[7\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_12385_ clknet_leaf_47_clk _01079_ VGND VGND VPWR VPWR data_array.data0\[14\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_10_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14124_ clknet_leaf_85_clk _02753_ VGND VGND VPWR VPWR data_array.data0\[1\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11336_ net950 net2620 net804 VGND VGND VPWR VPWR _03079_ sky130_fd_sc_hd__mux2_1
XFILLER_125_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14055_ clknet_leaf_37_clk _02684_ VGND VGND VPWR VPWR data_array.data1\[6\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_11267_ net962 net3653 net677 VGND VGND VPWR VPWR _03010_ sky130_fd_sc_hd__mux2_1
X_13006_ clknet_leaf_226_clk _01700_ VGND VGND VPWR VPWR data_array.data0\[3\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_10218_ net932 net4302 net360 VGND VGND VPWR VPWR _01965_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11198_ net981 net4296 net648 VGND VGND VPWR VPWR _02941_ sky130_fd_sc_hd__mux2_1
X_10149_ net949 net3264 net368 VGND VGND VPWR VPWR _01897_ sky130_fd_sc_hd__mux2_1
XFILLER_95_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13908_ clknet_leaf_86_clk _02537_ VGND VGND VPWR VPWR data_array.data1\[4\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_05690_ net19 fsm.tag_out0\[19\] VGND VGND VPWR VPWR _03207_ sky130_fd_sc_hd__and2b_1
XFILLER_36_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13839_ clknet_leaf_83_clk _02468_ VGND VGND VPWR VPWR data_array.data1\[3\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07360_ data_array.data0\[0\]\[56\] net1342 net1248 data_array.data0\[3\]\[56\] _04608_
+ VGND VGND VPWR VPWR _04609_ sky130_fd_sc_hd__a221o_1
X_06311_ tag_array.tag0\[0\]\[11\] net1401 net1307 tag_array.tag0\[3\]\[11\] _03654_
+ VGND VGND VPWR VPWR _03655_ sky130_fd_sc_hd__a221o_1
XFILLER_175_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07291_ data_array.data0\[13\]\[50\] net1537 net1441 data_array.data0\[14\]\[50\]
+ VGND VGND VPWR VPWR _04546_ sky130_fd_sc_hd__a22o_1
XFILLER_30_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09030_ net1839 net904 net418 VGND VGND VPWR VPWR _00785_ sky130_fd_sc_hd__mux2_1
XFILLER_50_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06242_ tag_array.tag0\[13\]\[5\] net1599 net1503 tag_array.tag0\[14\]\[5\] VGND
+ VGND VPWR VPWR _03592_ sky130_fd_sc_hd__a22o_1
XFILLER_164_829 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06173_ net1637 _03517_ net1211 _03525_ VGND VGND VPWR VPWR _03530_ sky130_fd_sc_hd__a22o_1
Xhold302 data_array.data0\[2\]\[23\] VGND VGND VPWR VPWR net1953 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold313 tag_array.dirty1\[1\] VGND VGND VPWR VPWR net1964 sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 data_array.data1\[4\]\[40\] VGND VGND VPWR VPWR net1975 sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 data_array.data1\[4\]\[37\] VGND VGND VPWR VPWR net1986 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold346 data_array.data0\[0\]\[14\] VGND VGND VPWR VPWR net1997 sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 data_array.data1\[2\]\[1\] VGND VGND VPWR VPWR net2008 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold368 data_array.data0\[1\]\[32\] VGND VGND VPWR VPWR net2019 sky130_fd_sc_hd__dlygate4sd3_1
X_09932_ net1102 net4123 net373 VGND VGND VPWR VPWR _01681_ sky130_fd_sc_hd__mux2_1
Xhold379 data_array.data1\[8\]\[37\] VGND VGND VPWR VPWR net2030 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout804 net805 VGND VGND VPWR VPWR net804 sky130_fd_sc_hd__buf_4
Xfanout815 _05360_ VGND VGND VPWR VPWR net815 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_74_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout837 net838 VGND VGND VPWR VPWR net837 sky130_fd_sc_hd__buf_6
X_09863_ net1019 net4467 net380 VGND VGND VPWR VPWR _01613_ sky130_fd_sc_hd__mux2_1
XFILLER_86_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout848 net849 VGND VGND VPWR VPWR net848 sky130_fd_sc_hd__buf_6
Xfanout859 _05546_ VGND VGND VPWR VPWR net859 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_98_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08814_ net2242 net989 net447 VGND VGND VPWR VPWR _00572_ sky130_fd_sc_hd__mux2_1
Xhold1002 tag_array.tag1\[9\]\[8\] VGND VGND VPWR VPWR net2653 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1013 data_array.data1\[9\]\[47\] VGND VGND VPWR VPWR net2664 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09794_ net1033 net2459 net391 VGND VGND VPWR VPWR _01545_ sky130_fd_sc_hd__mux2_1
Xhold1024 data_array.data0\[13\]\[9\] VGND VGND VPWR VPWR net2675 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1035 tag_array.tag1\[5\]\[11\] VGND VGND VPWR VPWR net2686 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1046 data_array.data1\[5\]\[52\] VGND VGND VPWR VPWR net2697 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1057 data_array.data1\[8\]\[2\] VGND VGND VPWR VPWR net2708 sky130_fd_sc_hd__dlygate4sd3_1
X_08745_ net743 net3954 net458 VGND VGND VPWR VPWR _00504_ sky130_fd_sc_hd__mux2_1
X_05957_ data_array.rdata0\[42\] net1666 net1148 VGND VGND VPWR VPWR _03432_ sky130_fd_sc_hd__o21a_1
Xhold1068 tag_array.tag1\[1\]\[23\] VGND VGND VPWR VPWR net2719 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1079 data_array.data0\[1\]\[27\] VGND VGND VPWR VPWR net2730 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08676_ net718 net2284 net494 VGND VGND VPWR VPWR _00435_ sky130_fd_sc_hd__mux2_1
X_05888_ data_array.rdata0\[19\] net850 net1147 VGND VGND VPWR VPWR _03386_ sky130_fd_sc_hd__o21a_1
XFILLER_26_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07627_ _04850_ _04851_ VGND VGND VPWR VPWR _00071_ sky130_fd_sc_hd__or2_1
XFILLER_53_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07558_ data_array.data1\[0\]\[10\] net1414 net1320 data_array.data1\[3\]\[10\] _04788_
+ VGND VGND VPWR VPWR _04789_ sky130_fd_sc_hd__a221o_1
XFILLER_167_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_157_3372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_472 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06509_ tag_array.tag1\[0\]\[4\] net1362 net1268 tag_array.tag1\[3\]\[4\] _03834_
+ VGND VGND VPWR VPWR _03835_ sky130_fd_sc_hd__a221o_1
X_07489_ data_array.data1\[13\]\[4\] net1584 net1488 data_array.data1\[14\]\[4\] VGND
+ VGND VPWR VPWR _04726_ sky130_fd_sc_hd__a22o_1
XFILLER_167_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_118_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09228_ net769 net2570 net647 VGND VGND VPWR VPWR _00982_ sky130_fd_sc_hd__mux2_1
XFILLER_6_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Left_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09159_ net907 net4077 net566 VGND VGND VPWR VPWR _00913_ sky130_fd_sc_hd__mux2_1
XFILLER_181_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12170_ clknet_leaf_170_clk _00978_ VGND VGND VPWR VPWR tag_array.tag0\[14\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11121_ net1035 net3369 net549 VGND VGND VPWR VPWR _02864_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_131_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold880 data_array.data0\[5\]\[11\] VGND VGND VPWR VPWR net2531 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold891 data_array.data0\[3\]\[42\] VGND VGND VPWR VPWR net2542 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11052_ net3159 net1052 net334 VGND VGND VPWR VPWR _02795_ sky130_fd_sc_hd__mux2_1
XFILLER_150_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10003_ net1074 net3978 net562 VGND VGND VPWR VPWR _01752_ sky130_fd_sc_hd__mux2_1
XFILLER_27_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2270 data_array.data0\[11\]\[33\] VGND VGND VPWR VPWR net3921 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2281 data_array.data0\[3\]\[39\] VGND VGND VPWR VPWR net3932 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2292 data_array.data0\[11\]\[0\] VGND VGND VPWR VPWR net3943 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1580 tag_array.tag1\[5\]\[7\] VGND VGND VPWR VPWR net3231 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1591 tag_array.tag1\[7\]\[8\] VGND VGND VPWR VPWR net3242 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_28_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11954_ clknet_leaf_30_clk _00762_ VGND VGND VPWR VPWR data_array.data0\[4\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10905_ net864 net4600 net517 VGND VGND VPWR VPWR _02650_ sky130_fd_sc_hd__mux2_1
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_177_3759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_192_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_192_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11885_ clknet_leaf_175_clk _00693_ VGND VGND VPWR VPWR data_array.data0\[5\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13624_ clknet_leaf_61_clk _02253_ VGND VGND VPWR VPWR data_array.data0\[9\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_177_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10836_ net1828 net886 net503 VGND VGND VPWR VPWR _02581_ sky130_fd_sc_hd__mux2_1
XFILLER_158_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13555_ clknet_leaf_212_clk _02184_ VGND VGND VPWR VPWR data_array.data1\[0\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10767_ net906 net2922 net490 VGND VGND VPWR VPWR _02512_ sky130_fd_sc_hd__mux2_1
XFILLER_34_1059 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12506_ clknet_leaf_203_clk _01200_ VGND VGND VPWR VPWR data_array.data1\[9\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13486_ clknet_leaf_159_clk _02116_ VGND VGND VPWR VPWR tag_array.tag0\[15\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_10698_ net3421 net924 net478 VGND VGND VPWR VPWR _02443_ sky130_fd_sc_hd__mux2_1
XFILLER_9_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12437_ clknet_leaf_16_clk _01131_ VGND VGND VPWR VPWR data_array.data0\[14\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_126_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12368_ clknet_leaf_256_clk _00045_ VGND VGND VPWR VPWR data_array.rdata0\[50\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_39_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14107_ clknet_leaf_60_clk _02736_ VGND VGND VPWR VPWR data_array.data0\[1\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_11319_ net1016 net2332 net798 VGND VGND VPWR VPWR _03062_ sky130_fd_sc_hd__mux2_1
XFILLER_113_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12299_ clknet_leaf_195_clk _01057_ VGND VGND VPWR VPWR tag_array.tag1\[12\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_56_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14038_ clknet_leaf_50_clk _02667_ VGND VGND VPWR VPWR data_array.data1\[6\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_141_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06860_ data_array.data0\[1\]\[11\] net1568 net1472 data_array.data0\[2\]\[11\] VGND
+ VGND VPWR VPWR _04154_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05811_ _03135_ fsm.tag_out0\[1\] _03170_ net1652 _03196_ VGND VGND VPWR VPWR _03328_
+ sky130_fd_sc_hd__a2111o_1
XFILLER_83_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06791_ _04090_ _04091_ VGND VGND VPWR VPWR _00044_ sky130_fd_sc_hd__or2_1
XFILLER_95_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08530_ net814 _05590_ net1700 VGND VGND VPWR VPWR _00304_ sky130_fd_sc_hd__a21o_1
X_05742_ net13 fsm.tag_out1\[13\] VGND VGND VPWR VPWR _03259_ sky130_fd_sc_hd__and2b_1
XFILLER_35_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08461_ net1129 _05543_ VGND VGND VPWR VPWR _05544_ sky130_fd_sc_hd__and2_1
XFILLER_36_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05673_ fsm.tag_out0\[14\] net14 VGND VGND VPWR VPWR _03190_ sky130_fd_sc_hd__and2b_1
XFILLER_35_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_183_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_183_clk
+ sky130_fd_sc_hd__clkbuf_8
X_07412_ data_array.data0\[9\]\[61\] net1553 net1457 data_array.data0\[10\]\[61\]
+ VGND VGND VPWR VPWR _04656_ sky130_fd_sc_hd__a22o_1
X_08392_ net1125 _05497_ VGND VGND VPWR VPWR _05498_ sky130_fd_sc_hd__and2_1
XFILLER_177_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07343_ data_array.data0\[12\]\[55\] net1343 net1249 data_array.data0\[15\]\[55\]
+ _04592_ VGND VGND VPWR VPWR _04593_ sky130_fd_sc_hd__a221o_1
XFILLER_32_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07274_ net1179 _04525_ _04529_ net1227 VGND VGND VPWR VPWR _04531_ sky130_fd_sc_hd__a22o_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09013_ net2328 net972 net419 VGND VGND VPWR VPWR _00768_ sky130_fd_sc_hd__mux2_1
X_06225_ tag_array.tag0\[8\]\[3\] net1373 net1280 tag_array.tag0\[11\]\[3\] _03576_
+ VGND VGND VPWR VPWR _03577_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_152_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold110 data_array.data0\[8\]\[15\] VGND VGND VPWR VPWR net1761 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06156_ net26 net27 VGND VGND VPWR VPWR _03513_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_76_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold121 data_array.data0\[8\]\[9\] VGND VGND VPWR VPWR net1772 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_160_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold132 data_array.data0\[2\]\[21\] VGND VGND VPWR VPWR net1783 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold143 tag_array.tag1\[1\]\[8\] VGND VGND VPWR VPWR net1794 sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 data_array.data0\[1\]\[51\] VGND VGND VPWR VPWR net1805 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 tag_array.tag1\[8\]\[8\] VGND VGND VPWR VPWR net1816 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_176_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06087_ data_array.rdata0\[2\] net1134 net1113 data_array.rdata1\[2\] VGND VGND VPWR
+ VPWR net285 sky130_fd_sc_hd__a22o_1
Xhold176 tag_array.tag1\[4\]\[18\] VGND VGND VPWR VPWR net1827 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold187 data_array.data1\[4\]\[23\] VGND VGND VPWR VPWR net1838 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout601 _05585_ VGND VGND VPWR VPWR net601 sky130_fd_sc_hd__buf_4
Xhold198 data_array.data1\[2\]\[22\] VGND VGND VPWR VPWR net1849 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout612 net614 VGND VGND VPWR VPWR net612 sky130_fd_sc_hd__buf_4
XFILLER_144_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09915_ net749 net4194 net602 VGND VGND VPWR VPWR _01665_ sky130_fd_sc_hd__mux2_1
XFILLER_99_982 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout623 _05567_ VGND VGND VPWR VPWR net623 sky130_fd_sc_hd__buf_2
XFILLER_132_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout634 net636 VGND VGND VPWR VPWR net634 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout645 net647 VGND VGND VPWR VPWR net645 sky130_fd_sc_hd__buf_4
Xfanout656 net660 VGND VGND VPWR VPWR net656 sky130_fd_sc_hd__clkbuf_8
X_09846_ net1085 net3865 net378 VGND VGND VPWR VPWR _01596_ sky130_fd_sc_hd__mux2_1
Xfanout667 net670 VGND VGND VPWR VPWR net667 sky130_fd_sc_hd__clkbuf_8
XFILLER_86_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout678 net679 VGND VGND VPWR VPWR net678 sky130_fd_sc_hd__buf_2
Xfanout689 net690 VGND VGND VPWR VPWR net689 sky130_fd_sc_hd__clkbuf_4
XFILLER_101_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09777_ net1102 net3241 net388 VGND VGND VPWR VPWR _01528_ sky130_fd_sc_hd__mux2_1
X_06989_ _04270_ _04271_ VGND VGND VPWR VPWR _00014_ sky130_fd_sc_hd__or2_1
XFILLER_37_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08728_ net2272 net710 net468 VGND VGND VPWR VPWR _00487_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_159_3412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_159_3423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08659_ net787 net3777 net496 VGND VGND VPWR VPWR _00418_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_174_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_174_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_15_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11670_ clknet_leaf_33_clk _00478_ VGND VGND VPWR VPWR tag_array.tag1\[1\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10621_ net2662 net977 net472 VGND VGND VPWR VPWR _02366_ sky130_fd_sc_hd__mux2_1
XFILLER_10_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_172_3667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13340_ clknet_leaf_53_clk _01970_ VGND VGND VPWR VPWR data_array.data0\[10\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
X_10552_ net997 net4583 net456 VGND VGND VPWR VPWR _02297_ sky130_fd_sc_hd__mux2_1
XFILLER_128_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13271_ clknet_leaf_84_clk _01901_ VGND VGND VPWR VPWR data_array.data0\[11\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10483_ net1012 net2554 net348 VGND VGND VPWR VPWR _02228_ sky130_fd_sc_hd__mux2_1
X_12222_ clknet_leaf_182_clk _00175_ VGND VGND VPWR VPWR fsm.tag_out1\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_142_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12153_ clknet_leaf_107_clk _00961_ VGND VGND VPWR VPWR tag_array.tag0\[13\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_97_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11104_ net1101 net2659 net542 VGND VGND VPWR VPWR _02847_ sky130_fd_sc_hd__mux2_1
XFILLER_151_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12084_ clknet_leaf_67_clk _00892_ VGND VGND VPWR VPWR data_array.data1\[14\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_111_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11035_ net1874 net860 net343 VGND VGND VPWR VPWR _02779_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_34_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_816 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12986_ clknet_leaf_262_clk _01680_ VGND VGND VPWR VPWR data_array.data0\[3\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11937_ clknet_leaf_45_clk _00745_ VGND VGND VPWR VPWR data_array.data0\[4\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_165_clk clknet_5_25__leaf_clk VGND VGND VPWR VPWR clknet_leaf_165_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_178_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11868_ clknet_leaf_270_clk _00676_ VGND VGND VPWR VPWR data_array.data0\[5\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_13607_ clknet_leaf_261_clk _02236_ VGND VGND VPWR VPWR data_array.data0\[9\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
X_10819_ net2022 net952 net503 VGND VGND VPWR VPWR _02564_ sky130_fd_sc_hd__mux2_1
XFILLER_60_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11799_ clknet_leaf_262_clk _00607_ VGND VGND VPWR VPWR data_array.data0\[7\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_158_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13538_ clknet_leaf_256_clk _02167_ VGND VGND VPWR VPWR data_array.data1\[0\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_146_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13469_ clknet_leaf_159_clk _02099_ VGND VGND VPWR VPWR tag_array.tag0\[15\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_174_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06010_ net153 net1156 _03466_ _03467_ VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__a22o_1
Xoutput204 net204 VGND VGND VPWR VPWR cpu_rdata[45] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_93_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput215 net215 VGND VGND VPWR VPWR cpu_rdata[55] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_93_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput226 net226 VGND VGND VPWR VPWR cpu_rdata[7] sky130_fd_sc_hd__buf_2
XFILLER_160_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput237 net237 VGND VGND VPWR VPWR mem_addr[16] sky130_fd_sc_hd__buf_2
XFILLER_153_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput248 net248 VGND VGND VPWR VPWR mem_addr[26] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput259 net259 VGND VGND VPWR VPWR mem_addr[7] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07961_ data_array.data1\[4\]\[47\] net1397 net1303 data_array.data1\[7\]\[47\] _05154_
+ VGND VGND VPWR VPWR _05155_ sky130_fd_sc_hd__a221o_1
XFILLER_141_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09700_ net789 net3211 net609 VGND VGND VPWR VPWR _01452_ sky130_fd_sc_hd__mux2_1
XFILLER_141_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06912_ _04200_ _04201_ VGND VGND VPWR VPWR _00006_ sky130_fd_sc_hd__or2_1
X_07892_ data_array.data1\[9\]\[41\] net1526 net1430 data_array.data1\[10\]\[41\]
+ VGND VGND VPWR VPWR _05092_ sky130_fd_sc_hd__a22o_1
XFILLER_114_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09631_ net762 net4426 net617 VGND VGND VPWR VPWR _01383_ sky130_fd_sc_hd__mux2_1
XFILLER_83_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06843_ data_array.data0\[0\]\[9\] net1389 net1295 data_array.data0\[3\]\[9\] _04138_
+ VGND VGND VPWR VPWR _04139_ sky130_fd_sc_hd__a221o_1
XFILLER_28_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09562_ net1102 net2819 net396 VGND VGND VPWR VPWR _01314_ sky130_fd_sc_hd__mux2_1
X_06774_ data_array.data0\[9\]\[3\] net1567 net1471 data_array.data0\[10\]\[3\] VGND
+ VGND VPWR VPWR _04076_ sky130_fd_sc_hd__a22o_1
XFILLER_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08513_ net1710 net607 VGND VGND VPWR VPWR _00299_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_19_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05725_ net10 fsm.tag_out1\[11\] VGND VGND VPWR VPWR _03242_ sky130_fd_sc_hd__xnor2_1
X_09493_ net755 net3878 net625 VGND VGND VPWR VPWR _01246_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_156_clk clknet_5_28__leaf_clk VGND VGND VPWR VPWR clknet_leaf_156_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_91_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08444_ net2255 net884 net687 VGND VGND VPWR VPWR _00277_ sky130_fd_sc_hd__mux2_1
X_05656_ fsm.tag_out0\[11\] net10 VGND VGND VPWR VPWR _03173_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_137_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08375_ net2348 net977 net691 VGND VGND VPWR VPWR _00254_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_154_3331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07326_ data_array.data0\[5\]\[53\] net1522 net1426 data_array.data0\[6\]\[53\] VGND
+ VGND VPWR VPWR _04578_ sky130_fd_sc_hd__a22o_1
XFILLER_165_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_150_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07257_ data_array.data0\[4\]\[47\] net1387 net1293 data_array.data0\[7\]\[47\] _04514_
+ VGND VGND VPWR VPWR _04515_ sky130_fd_sc_hd__a221o_1
XFILLER_164_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06208_ _03560_ _03561_ VGND VGND VPWR VPWR _00142_ sky130_fd_sc_hd__or2_1
XFILLER_124_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07188_ data_array.data0\[9\]\[41\] net1527 net1431 data_array.data0\[10\]\[41\]
+ VGND VGND VPWR VPWR _04452_ sky130_fd_sc_hd__a22o_1
XFILLER_180_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06139_ data_array.rdata0\[54\] net1136 net1117 data_array.rdata1\[54\] VGND VGND
+ VPWR VPWR net312 sky130_fd_sc_hd__a22o_1
XFILLER_160_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1407 net1408 VGND VGND VPWR VPWR net1407 sky130_fd_sc_hd__clkbuf_4
XFILLER_105_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout420 net421 VGND VGND VPWR VPWR net420 sky130_fd_sc_hd__buf_4
XFILLER_63_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1418 net1421 VGND VGND VPWR VPWR net1418 sky130_fd_sc_hd__clkbuf_4
Xfanout431 net433 VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__buf_4
Xfanout1429 net1430 VGND VGND VPWR VPWR net1429 sky130_fd_sc_hd__clkbuf_4
XFILLER_87_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout442 net443 VGND VGND VPWR VPWR net442 sky130_fd_sc_hd__buf_4
Xfanout453 net459 VGND VGND VPWR VPWR net453 sky130_fd_sc_hd__buf_4
Xfanout464 net465 VGND VGND VPWR VPWR net464 sky130_fd_sc_hd__clkbuf_4
Xfanout475 net476 VGND VGND VPWR VPWR net475 sky130_fd_sc_hd__buf_4
Xfanout486 net489 VGND VGND VPWR VPWR net486 sky130_fd_sc_hd__buf_4
XFILLER_171_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout497 net499 VGND VGND VPWR VPWR net497 sky130_fd_sc_hd__buf_4
X_09829_ net894 net4087 net388 VGND VGND VPWR VPWR _01580_ sky130_fd_sc_hd__mux2_1
XFILLER_150_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1069 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12840_ clknet_leaf_17_clk _01534_ VGND VGND VPWR VPWR data_array.data0\[12\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_126_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ clknet_leaf_173_clk _01465_ VGND VGND VPWR VPWR tag_array.tag0\[6\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_147_clk clknet_5_31__leaf_clk VGND VGND VPWR VPWR clknet_leaf_147_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_174_3707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ clknet_leaf_137_clk _00530_ VGND VGND VPWR VPWR tag_array.tag0\[9\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_727 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14441_ clknet_leaf_267_clk _03064_ VGND VGND VPWR VPWR data_array.data1\[7\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_11653_ clknet_leaf_100_clk _00461_ VGND VGND VPWR VPWR tag_array.tag1\[2\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_10604_ net2304 net1044 net469 VGND VGND VPWR VPWR _02349_ sky130_fd_sc_hd__mux2_1
XFILLER_156_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14372_ clknet_leaf_24_clk _02995_ VGND VGND VPWR VPWR data_array.data1\[10\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11584_ clknet_leaf_97_clk _00392_ VGND VGND VPWR VPWR tag_array.tag1\[4\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_168_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13323_ clknet_leaf_261_clk _01953_ VGND VGND VPWR VPWR data_array.data0\[10\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10535_ net1066 net3352 net460 VGND VGND VPWR VPWR _02280_ sky130_fd_sc_hd__mux2_1
XFILLER_13_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13254_ clknet_leaf_229_clk _01884_ VGND VGND VPWR VPWR data_array.data0\[11\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10466_ net1081 net3707 net350 VGND VGND VPWR VPWR _02211_ sky130_fd_sc_hd__mux2_1
XFILLER_89_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12205_ clknet_leaf_153_clk _00134_ VGND VGND VPWR VPWR fsm.tag_out0\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_142_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13185_ clknet_leaf_12_clk _00078_ VGND VGND VPWR VPWR data_array.rdata1\[22\] sky130_fd_sc_hd__dfxtp_1
X_10397_ net2192 net1067 net667 VGND VGND VPWR VPWR _02143_ sky130_fd_sc_hd__mux2_1
XFILLER_69_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12136_ clknet_leaf_181_clk _00944_ VGND VGND VPWR VPWR tag_array.tag0\[12\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_123_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_941 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12067_ clknet_leaf_200_clk _00875_ VGND VGND VPWR VPWR data_array.data1\[14\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_111_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Left_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11018_ net2136 net928 net337 VGND VGND VPWR VPWR _02762_ sky130_fd_sc_hd__mux2_1
XFILLER_37_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1070 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_138_clk clknet_5_31__leaf_clk VGND VGND VPWR VPWR clknet_leaf_138_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12969_ clknet_leaf_160_clk _01663_ VGND VGND VPWR VPWR tag_array.tag0\[4\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06490_ tag_array.tag1\[1\]\[2\] net1541 net1445 tag_array.tag1\[2\]\[2\] VGND VGND
+ VPWR VPWR _03818_ sky130_fd_sc_hd__a22o_1
XFILLER_178_537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08160_ tag_array.dirty0\[9\] net1593 net1497 tag_array.dirty0\[10\] VGND VGND VPWR
+ VPWR _05336_ sky130_fd_sc_hd__a22o_1
XFILLER_158_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07111_ data_array.data0\[13\]\[34\] net1531 net1435 data_array.data0\[14\]\[34\]
+ VGND VGND VPWR VPWR _04382_ sky130_fd_sc_hd__a22o_1
XFILLER_118_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08091_ data_array.data1\[8\]\[59\] net1381 net1287 data_array.data1\[11\]\[59\]
+ _05272_ VGND VGND VPWR VPWR _05273_ sky130_fd_sc_hd__a221o_1
XFILLER_174_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload30 clknet_leaf_10_clk VGND VGND VPWR VPWR clkload30/Y sky130_fd_sc_hd__clkinv_4
XFILLER_146_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07042_ net1619 _04313_ _04317_ net1193 VGND VGND VPWR VPWR _04320_ sky130_fd_sc_hd__a22o_1
Xclkload41 clknet_leaf_21_clk VGND VGND VPWR VPWR clkload41/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_106_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload52 clknet_leaf_250_clk VGND VGND VPWR VPWR clkload52/Y sky130_fd_sc_hd__inv_6
Xclkload63 clknet_leaf_241_clk VGND VGND VPWR VPWR clkload63/Y sky130_fd_sc_hd__bufinv_16
XFILLER_161_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload74 clknet_leaf_240_clk VGND VGND VPWR VPWR clkload74/Y sky130_fd_sc_hd__clkinv_2
XFILLER_47_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload85 clknet_leaf_45_clk VGND VGND VPWR VPWR clkload85/X sky130_fd_sc_hd__clkbuf_4
Xclkload96 clknet_leaf_58_clk VGND VGND VPWR VPWR clkload96/Y sky130_fd_sc_hd__inv_8
XFILLER_47_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08993_ net1977 net1052 net423 VGND VGND VPWR VPWR _00748_ sky130_fd_sc_hd__mux2_1
Xhold2803 data_array.data1\[11\]\[28\] VGND VGND VPWR VPWR net4454 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_173_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2814 tag_array.tag1\[11\]\[19\] VGND VGND VPWR VPWR net4465 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2825 tag_array.tag0\[9\]\[16\] VGND VGND VPWR VPWR net4476 sky130_fd_sc_hd__dlygate4sd3_1
X_07944_ net1192 _05133_ _05137_ net1618 VGND VGND VPWR VPWR _05140_ sky130_fd_sc_hd__a22o_1
Xhold2836 data_array.data1\[6\]\[32\] VGND VGND VPWR VPWR net4487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2847 data_array.data0\[11\]\[32\] VGND VGND VPWR VPWR net4498 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2858 data_array.data1\[14\]\[48\] VGND VGND VPWR VPWR net4509 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_147_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2869 tag_array.tag0\[0\]\[16\] VGND VGND VPWR VPWR net4520 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07875_ data_array.data1\[12\]\[39\] net1347 net1253 data_array.data1\[15\]\[39\]
+ _05076_ VGND VGND VPWR VPWR _05077_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_3_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09614_ net894 net3654 net396 VGND VGND VPWR VPWR _01366_ sky130_fd_sc_hd__mux2_1
X_06826_ data_array.data0\[12\]\[8\] net1343 net1249 data_array.data0\[15\]\[8\] _04122_
+ VGND VGND VPWR VPWR _04123_ sky130_fd_sc_hd__a221o_1
X_09545_ net748 net4335 net619 VGND VGND VPWR VPWR _01298_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_129_clk clknet_5_30__leaf_clk VGND VGND VPWR VPWR clknet_leaf_129_clk
+ sky130_fd_sc_hd__clkbuf_8
X_06757_ net1213 _04055_ _04059_ net1165 VGND VGND VPWR VPWR _04061_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_174_Right_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05708_ _03194_ _03196_ _03199_ _03224_ VGND VGND VPWR VPWR _03225_ sky130_fd_sc_hd__or4_1
X_09476_ net725 net3526 net658 VGND VGND VPWR VPWR _01229_ sky130_fd_sc_hd__mux2_1
X_06688_ tag_array.tag1\[5\]\[20\] net1541 net1445 tag_array.tag1\[6\]\[20\] VGND
+ VGND VPWR VPWR _03998_ sky130_fd_sc_hd__a22o_1
XFILLER_51_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08427_ net145 net80 net1638 VGND VGND VPWR VPWR _05521_ sky130_fd_sc_hd__mux2_1
XFILLER_24_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05639_ net25 fsm.tag_out0\[24\] VGND VGND VPWR VPWR _03156_ sky130_fd_sc_hd__xor2_1
XFILLER_138_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08358_ net119 net54 net1638 VGND VGND VPWR VPWR _05475_ sky130_fd_sc_hd__mux2_1
Xclkload2 clknet_5_4__leaf_clk VGND VGND VPWR VPWR clkload2/Y sky130_fd_sc_hd__inv_6
X_07309_ data_array.data0\[13\]\[52\] net1549 net1453 data_array.data0\[14\]\[52\]
+ VGND VGND VPWR VPWR _04562_ sky130_fd_sc_hd__a22o_1
XFILLER_149_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08289_ net154 net89 net1643 VGND VGND VPWR VPWR _05429_ sky130_fd_sc_hd__mux2_1
XFILLER_125_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10320_ net3870 net882 net636 VGND VGND VPWR VPWR _02067_ sky130_fd_sc_hd__mux2_1
XFILLER_180_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10251_ net739 net3447 net597 VGND VGND VPWR VPWR _01998_ sky130_fd_sc_hd__mux2_1
XFILLER_152_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_167_3566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10182_ net1077 net3684 net355 VGND VGND VPWR VPWR _01929_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_167_3577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1204 net1206 VGND VGND VPWR VPWR net1204 sky130_fd_sc_hd__buf_4
Xfanout1215 net1223 VGND VGND VPWR VPWR net1215 sky130_fd_sc_hd__clkbuf_4
Xfanout1226 net1228 VGND VGND VPWR VPWR net1226 sky130_fd_sc_hd__buf_4
Xfanout1237 net1282 VGND VGND VPWR VPWR net1237 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_184_3891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1248 net1258 VGND VGND VPWR VPWR net1248 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_128_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1259 net1261 VGND VGND VPWR VPWR net1259 sky130_fd_sc_hd__clkbuf_4
XFILLER_75_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13941_ clknet_leaf_25_clk _02570_ VGND VGND VPWR VPWR data_array.data1\[4\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
X_13872_ clknet_leaf_123_clk _02501_ VGND VGND VPWR VPWR data_array.data1\[3\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_87 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12823_ clknet_leaf_140_clk _01517_ VGND VGND VPWR VPWR tag_array.tag1\[0\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_141_Right_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12754_ clknet_leaf_178_clk _01448_ VGND VGND VPWR VPWR tag_array.tag0\[5\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11705_ clknet_leaf_100_clk _00513_ VGND VGND VPWR VPWR tag_array.tag1\[15\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12685_ clknet_leaf_179_clk _01379_ VGND VGND VPWR VPWR tag_array.tag0\[8\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_14424_ clknet_leaf_28_clk _03047_ VGND VGND VPWR VPWR data_array.data1\[7\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_11636_ clknet_leaf_31_clk _00444_ VGND VGND VPWR VPWR tag_array.tag1\[2\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_128_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11567_ clknet_leaf_141_clk _00375_ VGND VGND VPWR VPWR tag_array.tag1\[5\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_14355_ clknet_leaf_199_clk _02978_ VGND VGND VPWR VPWR data_array.data1\[10\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13306_ clknet_leaf_63_clk _01936_ VGND VGND VPWR VPWR data_array.data0\[10\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_155_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10518_ net873 net3644 net348 VGND VGND VPWR VPWR _02263_ sky130_fd_sc_hd__mux2_1
X_14286_ clknet_leaf_268_clk _02915_ VGND VGND VPWR VPWR data_array.data1\[11\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold709 tag_array.tag0\[6\]\[16\] VGND VGND VPWR VPWR net2360 sky130_fd_sc_hd__dlygate4sd3_1
X_11498_ clknet_leaf_172_clk _00306_ VGND VGND VPWR VPWR tag_array.valid1\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_90_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13237_ clknet_leaf_111_clk _01867_ VGND VGND VPWR VPWR data_array.data0\[11\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_10449_ net2271 net858 net664 VGND VGND VPWR VPWR _02195_ sky130_fd_sc_hd__mux2_1
XFILLER_130_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13168_ clknet_leaf_202_clk _00119_ VGND VGND VPWR VPWR data_array.rdata1\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_151_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12119_ clknet_leaf_163_clk _00927_ VGND VGND VPWR VPWR tag_array.tag0\[12\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_05990_ data_array.rdata0\[53\] net846 net1142 VGND VGND VPWR VPWR _03454_ sky130_fd_sc_hd__o21a_1
X_13099_ clknet_leaf_245_clk _01793_ VGND VGND VPWR VPWR data_array.data1\[13\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1409 tag_array.dirty0\[15\] VGND VGND VPWR VPWR net3060 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_88_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07660_ _04880_ _04881_ VGND VGND VPWR VPWR _00074_ sky130_fd_sc_hd__or2_1
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_914 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06611_ tag_array.tag1\[1\]\[13\] net1611 net1515 tag_array.tag1\[2\]\[13\] VGND
+ VGND VPWR VPWR _03928_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_49_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07591_ data_array.data1\[4\]\[13\] net1359 net1265 data_array.data1\[7\]\[13\] _04818_
+ VGND VGND VPWR VPWR _04819_ sky130_fd_sc_hd__a221o_1
X_09330_ net1080 net2948 net408 VGND VGND VPWR VPWR _01083_ sky130_fd_sc_hd__mux2_1
X_06542_ tag_array.tag1\[4\]\[7\] net1420 net1326 tag_array.tag1\[7\]\[7\] _03864_
+ VGND VGND VPWR VPWR _03865_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_66_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_857 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09261_ net734 net3605 net569 VGND VGND VPWR VPWR _01015_ sky130_fd_sc_hd__mux2_1
X_06473_ tag_array.tag1\[13\]\[1\] net1560 net1464 tag_array.tag1\[14\]\[1\] VGND
+ VGND VPWR VPWR _03802_ sky130_fd_sc_hd__a22o_1
X_08212_ net1649 net1158 net5 VGND VGND VPWR VPWR _05376_ sky130_fd_sc_hd__and3_1
X_09192_ net713 net2843 net627 VGND VGND VPWR VPWR _00946_ sky130_fd_sc_hd__mux2_1
XFILLER_140_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08143_ net1171 _05315_ _05319_ net1219 VGND VGND VPWR VPWR _05321_ sky130_fd_sc_hd__a22o_1
XFILLER_14_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08074_ data_array.data1\[5\]\[57\] net1528 net1432 data_array.data1\[6\]\[57\] VGND
+ VGND VPWR VPWR _05258_ sky130_fd_sc_hd__a22o_1
Xclkload130 clknet_leaf_86_clk VGND VGND VPWR VPWR clkload130/Y sky130_fd_sc_hd__clkinv_8
XFILLER_162_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload141 clknet_leaf_223_clk VGND VGND VPWR VPWR clkload141/Y sky130_fd_sc_hd__bufinv_16
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload152 clknet_leaf_229_clk VGND VGND VPWR VPWR clkload152/Y sky130_fd_sc_hd__inv_6
XFILLER_128_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload163 clknet_leaf_201_clk VGND VGND VPWR VPWR clkload163/X sky130_fd_sc_hd__clkbuf_8
XFILLER_134_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07025_ data_array.data0\[5\]\[26\] net1528 net1432 data_array.data0\[6\]\[26\] VGND
+ VGND VPWR VPWR _04304_ sky130_fd_sc_hd__a22o_1
Xclkload174 clknet_leaf_199_clk VGND VGND VPWR VPWR clkload174/Y sky130_fd_sc_hd__clkinv_4
Xclkload185 clknet_leaf_186_clk VGND VGND VPWR VPWR clkload185/Y sky130_fd_sc_hd__inv_6
Xclkload196 clknet_leaf_166_clk VGND VGND VPWR VPWR clkload196/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_149_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2600 tag_array.tag1\[12\]\[14\] VGND VGND VPWR VPWR net4251 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2611 data_array.data0\[15\]\[36\] VGND VGND VPWR VPWR net4262 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2622 data_array.data1\[15\]\[39\] VGND VGND VPWR VPWR net4273 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2633 data_array.data0\[14\]\[20\] VGND VGND VPWR VPWR net4284 sky130_fd_sc_hd__dlygate4sd3_1
X_08976_ net860 net3179 net433 VGND VGND VPWR VPWR _00732_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_145_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2644 data_array.data1\[15\]\[44\] VGND VGND VPWR VPWR net4295 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1910 data_array.data1\[13\]\[23\] VGND VGND VPWR VPWR net3561 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2655 data_array.data0\[12\]\[58\] VGND VGND VPWR VPWR net4306 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 tag_array.valid1\[5\] VGND VGND VPWR VPWR net1698 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07927_ data_array.data1\[1\]\[44\] net1589 net1493 data_array.data1\[2\]\[44\] VGND
+ VGND VPWR VPWR _05124_ sky130_fd_sc_hd__a22o_1
Xhold1921 data_array.data0\[15\]\[20\] VGND VGND VPWR VPWR net3572 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2666 data_array.data0\[15\]\[57\] VGND VGND VPWR VPWR net4317 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 tag_array.valid1\[15\] VGND VGND VPWR VPWR net1709 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1932 lru_array.lru_mem\[3\] VGND VGND VPWR VPWR net3583 sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 tag_array.valid0\[8\] VGND VGND VPWR VPWR net1720 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2677 data_array.data0\[13\]\[33\] VGND VGND VPWR VPWR net4328 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_162_3474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1943 data_array.data1\[5\]\[39\] VGND VGND VPWR VPWR net3594 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2688 data_array.data0\[7\]\[38\] VGND VGND VPWR VPWR net4339 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_162_3485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2699 tag_array.tag1\[15\]\[9\] VGND VGND VPWR VPWR net4350 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_21_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1954 tag_array.tag1\[14\]\[14\] VGND VGND VPWR VPWR net3605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1965 tag_array.tag0\[4\]\[12\] VGND VGND VPWR VPWR net3616 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07858_ _05060_ _05061_ VGND VGND VPWR VPWR _00094_ sky130_fd_sc_hd__or2_1
XFILLER_84_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1976 tag_array.tag0\[9\]\[11\] VGND VGND VPWR VPWR net3627 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1987 data_array.data0\[15\]\[48\] VGND VGND VPWR VPWR net3638 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1998 data_array.data1\[12\]\[38\] VGND VGND VPWR VPWR net3649 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_123_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06809_ data_array.data0\[5\]\[6\] net1521 net1425 data_array.data0\[6\]\[6\] VGND
+ VGND VPWR VPWR _04108_ sky130_fd_sc_hd__a22o_1
X_07789_ data_array.data1\[0\]\[31\] net1381 net1287 data_array.data1\[3\]\[31\] _04998_
+ VGND VGND VPWR VPWR _04999_ sky130_fd_sc_hd__a221o_1
X_09528_ net717 net4563 net622 VGND VGND VPWR VPWR _01281_ sky130_fd_sc_hd__mux2_1
X_09459_ net791 net2492 net655 VGND VGND VPWR VPWR _01212_ sky130_fd_sc_hd__mux2_1
XFILLER_101_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12470_ clknet_leaf_24_clk _01164_ VGND VGND VPWR VPWR data_array.data1\[9\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11421_ clknet_leaf_112_clk _00231_ VGND VGND VPWR VPWR data_array.data0\[0\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_138_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14140_ clknet_leaf_223_clk _02769_ VGND VGND VPWR VPWR data_array.data0\[1\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_3606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11352_ net886 net3416 net796 VGND VGND VPWR VPWR _03095_ sky130_fd_sc_hd__mux2_1
XFILLER_180_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_169_3617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10303_ net2288 net950 net642 VGND VGND VPWR VPWR _02050_ sky130_fd_sc_hd__mux2_1
X_14071_ clknet_leaf_74_clk _02700_ VGND VGND VPWR VPWR data_array.data1\[6\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_89_Left_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11283_ net899 net4314 net673 VGND VGND VPWR VPWR _03026_ sky130_fd_sc_hd__mux2_1
X_13022_ clknet_leaf_218_clk _01716_ VGND VGND VPWR VPWR data_array.data0\[3\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
X_10234_ net869 net3606 net361 VGND VGND VPWR VPWR _01981_ sky130_fd_sc_hd__mux2_1
Xfanout1001 _05474_ VGND VGND VPWR VPWR net1001 sky130_fd_sc_hd__buf_1
Xfanout1012 _05468_ VGND VGND VPWR VPWR net1012 sky130_fd_sc_hd__clkbuf_2
X_10165_ net884 net4526 net363 VGND VGND VPWR VPWR _01913_ sky130_fd_sc_hd__mux2_1
Xfanout1023 _05464_ VGND VGND VPWR VPWR net1023 sky130_fd_sc_hd__clkbuf_2
Xfanout1034 _05458_ VGND VGND VPWR VPWR net1034 sky130_fd_sc_hd__clkbuf_2
Xfanout1045 _05452_ VGND VGND VPWR VPWR net1045 sky130_fd_sc_hd__buf_1
Xfanout1056 _05446_ VGND VGND VPWR VPWR net1056 sky130_fd_sc_hd__clkbuf_2
XFILLER_121_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10096_ net1855 net741 net642 VGND VGND VPWR VPWR _01845_ sky130_fd_sc_hd__mux2_1
Xfanout1067 _05442_ VGND VGND VPWR VPWR net1067 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1078 net1079 VGND VGND VPWR VPWR net1078 sky130_fd_sc_hd__clkbuf_2
Xfanout1089 _05430_ VGND VGND VPWR VPWR net1089 sky130_fd_sc_hd__clkbuf_2
X_13924_ clknet_leaf_30_clk _02553_ VGND VGND VPWR VPWR data_array.data1\[4\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_98_Left_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13855_ clknet_leaf_200_clk _02484_ VGND VGND VPWR VPWR data_array.data1\[3\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12806_ clknet_leaf_188_clk _01500_ VGND VGND VPWR VPWR tag_array.tag1\[10\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_10998_ net1752 net1009 net336 VGND VGND VPWR VPWR _02742_ sky130_fd_sc_hd__mux2_1
X_13786_ clknet_leaf_18_clk _02415_ VGND VGND VPWR VPWR data_array.data1\[2\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_163_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1032 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ clknet_leaf_143_clk _01431_ VGND VGND VPWR VPWR tag_array.tag0\[5\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_26_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12668_ clknet_leaf_25_clk _01362_ VGND VGND VPWR VPWR data_array.data0\[15\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14407_ clknet_leaf_238_clk _03030_ VGND VGND VPWR VPWR data_array.data1\[10\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
X_11619_ clknet_leaf_102_clk _00427_ VGND VGND VPWR VPWR tag_array.tag1\[3\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_12599_ clknet_leaf_180_clk _01293_ VGND VGND VPWR VPWR tag_array.tag0\[0\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14338_ clknet_leaf_203_clk _02967_ VGND VGND VPWR VPWR data_array.data1\[11\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold506 data_array.data1\[6\]\[15\] VGND VGND VPWR VPWR net2157 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold517 data_array.data0\[2\]\[29\] VGND VGND VPWR VPWR net2168 sky130_fd_sc_hd__dlygate4sd3_1
Xhold528 tag_array.tag1\[8\]\[18\] VGND VGND VPWR VPWR net2179 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold539 data_array.data1\[0\]\[9\] VGND VGND VPWR VPWR net2190 sky130_fd_sc_hd__dlygate4sd3_1
X_14269_ clknet_leaf_5_clk _02898_ VGND VGND VPWR VPWR data_array.data1\[12\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_855 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08830_ net2250 net927 net442 VGND VGND VPWR VPWR _00588_ sky130_fd_sc_hd__mux2_1
XFILLER_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1206 tag_array.tag0\[15\]\[14\] VGND VGND VPWR VPWR net2857 sky130_fd_sc_hd__dlygate4sd3_1
X_08761_ net781 net4496 net450 VGND VGND VPWR VPWR _00520_ sky130_fd_sc_hd__mux2_1
XFILLER_100_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1217 tag_array.tag1\[0\]\[10\] VGND VGND VPWR VPWR net2868 sky130_fd_sc_hd__dlygate4sd3_1
X_05973_ data_array.rdata1\[47\] net833 net842 VGND VGND VPWR VPWR _03443_ sky130_fd_sc_hd__a21o_1
Xhold1228 tag_array.tag0\[15\]\[21\] VGND VGND VPWR VPWR net2879 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1239 data_array.data1\[12\]\[23\] VGND VGND VPWR VPWR net2890 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07712_ data_array.data1\[0\]\[24\] net1387 net1293 data_array.data1\[3\]\[24\] _04928_
+ VGND VGND VPWR VPWR _04929_ sky130_fd_sc_hd__a221o_1
Xfanout1590 net1591 VGND VGND VPWR VPWR net1590 sky130_fd_sc_hd__buf_2
X_08692_ net3032 net756 net487 VGND VGND VPWR VPWR _00451_ sky130_fd_sc_hd__mux2_1
XFILLER_26_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07643_ data_array.data1\[13\]\[18\] net1568 net1472 data_array.data1\[14\]\[18\]
+ VGND VGND VPWR VPWR _04866_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_140_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07574_ data_array.data1\[8\]\[12\] net1395 net1301 data_array.data1\[11\]\[12\]
+ _04802_ VGND VGND VPWR VPWR _04803_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_101_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09313_ net728 net2700 net551 VGND VGND VPWR VPWR _01067_ sky130_fd_sc_hd__mux2_1
X_06525_ net1636 _03843_ _03847_ net1210 VGND VGND VPWR VPWR _03850_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_81_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_310 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_60_clk clknet_5_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_60_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_21_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09244_ net704 net3445 net647 VGND VGND VPWR VPWR _00998_ sky130_fd_sc_hd__mux2_1
XFILLER_90_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06456_ tag_array.tag0\[12\]\[24\] net1374 net1281 tag_array.tag0\[15\]\[24\] _03786_
+ VGND VGND VPWR VPWR _03787_ sky130_fd_sc_hd__a221o_1
XFILLER_178_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09175_ net781 net3195 net627 VGND VGND VPWR VPWR _00929_ sky130_fd_sc_hd__mux2_1
X_06387_ tag_array.tag0\[1\]\[18\] net1564 net1468 tag_array.tag0\[2\]\[18\] VGND
+ VGND VPWR VPWR _03724_ sky130_fd_sc_hd__a22o_1
XFILLER_175_860 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08126_ data_array.data1\[4\]\[62\] net1415 net1321 data_array.data1\[7\]\[62\] _05304_
+ VGND VGND VPWR VPWR _05305_ sky130_fd_sc_hd__a221o_1
XFILLER_135_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08057_ data_array.data1\[13\]\[56\] net1532 net1436 data_array.data1\[14\]\[56\]
+ VGND VGND VPWR VPWR _05242_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_79_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07008_ data_array.data0\[0\]\[24\] net1386 net1292 data_array.data0\[3\]\[24\] _04288_
+ VGND VGND VPWR VPWR _04289_ sky130_fd_sc_hd__a221o_1
XFILLER_134_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput104 mem_rdata[14] VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_1
XFILLER_103_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput115 mem_rdata[24] VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_1
XFILLER_163_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput126 mem_rdata[34] VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_1
Xhold2430 data_array.data0\[10\]\[11\] VGND VGND VPWR VPWR net4081 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput137 mem_rdata[44] VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_1
Xhold2441 data_array.data0\[11\]\[24\] VGND VGND VPWR VPWR net4092 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2452 data_array.data1\[3\]\[16\] VGND VGND VPWR VPWR net4103 sky130_fd_sc_hd__dlygate4sd3_1
Xinput148 mem_rdata[54] VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_1
Xinput159 mem_rdata[6] VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_1
Xhold2463 data_array.data0\[7\]\[34\] VGND VGND VPWR VPWR net4114 sky130_fd_sc_hd__dlygate4sd3_1
X_08959_ net928 net2801 net427 VGND VGND VPWR VPWR _00715_ sky130_fd_sc_hd__mux2_1
Xhold2474 tag_array.tag1\[5\]\[5\] VGND VGND VPWR VPWR net4125 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_5_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2485 tag_array.dirty0\[8\] VGND VGND VPWR VPWR net4136 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1740 data_array.data0\[14\]\[29\] VGND VGND VPWR VPWR net3391 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1751 data_array.data1\[3\]\[23\] VGND VGND VPWR VPWR net3402 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2496 data_array.data0\[7\]\[39\] VGND VGND VPWR VPWR net4147 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1762 tag_array.tag0\[8\]\[14\] VGND VGND VPWR VPWR net3413 sky130_fd_sc_hd__dlygate4sd3_1
X_11970_ clknet_leaf_87_clk _00778_ VGND VGND VPWR VPWR data_array.data0\[4\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1773 data_array.data1\[14\]\[60\] VGND VGND VPWR VPWR net3424 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_5_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1784 tag_array.tag0\[3\]\[16\] VGND VGND VPWR VPWR net3435 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_179_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1795 data_array.data0\[5\]\[5\] VGND VGND VPWR VPWR net3446 sky130_fd_sc_hd__dlygate4sd3_1
X_10921_ net1056 net4141 net528 VGND VGND VPWR VPWR _02666_ sky130_fd_sc_hd__mux2_1
XFILLER_56_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13640_ clknet_leaf_226_clk _02269_ VGND VGND VPWR VPWR data_array.data1\[15\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_10852_ net1078 net2660 net519 VGND VGND VPWR VPWR _02597_ sky130_fd_sc_hd__mux2_1
XFILLER_32_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_179_3790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13571_ clknet_leaf_29_clk _02200_ VGND VGND VPWR VPWR tag_array.dirty1\[3\] sky130_fd_sc_hd__dfxtp_1
X_10783_ net2363 net1098 net507 VGND VGND VPWR VPWR _02528_ sky130_fd_sc_hd__mux2_1
XFILLER_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_51_clk clknet_5_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_51_clk sky130_fd_sc_hd__clkbuf_8
X_12522_ clknet_leaf_195_clk _01216_ VGND VGND VPWR VPWR tag_array.tag1\[11\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12453_ clknet_leaf_199_clk _01147_ VGND VGND VPWR VPWR data_array.data1\[9\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_11404_ clknet_leaf_189_clk _00214_ VGND VGND VPWR VPWR tag_array.tag1\[7\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12384_ clknet_leaf_247_clk _01078_ VGND VGND VPWR VPWR data_array.data0\[14\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_181_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14123_ clknet_leaf_244_clk _02752_ VGND VGND VPWR VPWR data_array.data0\[1\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
X_11335_ net952 net3905 net796 VGND VGND VPWR VPWR _03078_ sky130_fd_sc_hd__mux2_1
XFILLER_4_553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11266_ net966 net4309 net681 VGND VGND VPWR VPWR _03009_ sky130_fd_sc_hd__mux2_1
X_14054_ clknet_leaf_70_clk _02683_ VGND VGND VPWR VPWR data_array.data1\[6\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_13005_ clknet_leaf_125_clk _01699_ VGND VGND VPWR VPWR data_array.data0\[3\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_97_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10217_ net939 net3967 net358 VGND VGND VPWR VPWR _01964_ sky130_fd_sc_hd__mux2_1
XFILLER_97_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11197_ net984 net2899 net655 VGND VGND VPWR VPWR _02940_ sky130_fd_sc_hd__mux2_1
XFILLER_122_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10148_ net955 net4012 net369 VGND VGND VPWR VPWR _01896_ sky130_fd_sc_hd__mux2_1
XFILLER_48_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_85_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10079_ net708 net2080 net601 VGND VGND VPWR VPWR _01828_ sky130_fd_sc_hd__mux2_1
X_13907_ clknet_leaf_35_clk _02536_ VGND VGND VPWR VPWR data_array.data1\[4\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13838_ clknet_leaf_268_clk _02467_ VGND VGND VPWR VPWR data_array.data1\[3\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_63_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13769_ clknet_leaf_267_clk _02398_ VGND VGND VPWR VPWR data_array.data1\[2\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_42_clk clknet_5_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_42_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_31_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06310_ tag_array.tag0\[1\]\[11\] net1592 net1496 tag_array.tag0\[2\]\[11\] VGND
+ VGND VPWR VPWR _03654_ sky130_fd_sc_hd__a22o_1
XFILLER_148_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07290_ data_array.data0\[4\]\[50\] net1346 net1252 data_array.data0\[7\]\[50\] _04544_
+ VGND VGND VPWR VPWR _04545_ sky130_fd_sc_hd__a221o_1
XFILLER_31_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06241_ _03590_ _03591_ VGND VGND VPWR VPWR _00150_ sky130_fd_sc_hd__or2_1
XFILLER_148_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06172_ tag_array.valid0\[4\] net1407 net1313 tag_array.valid0\[7\] _03528_ VGND
+ VGND VPWR VPWR _03529_ sky130_fd_sc_hd__a221o_1
Xhold303 data_array.data1\[8\]\[59\] VGND VGND VPWR VPWR net1954 sky130_fd_sc_hd__dlygate4sd3_1
Xhold314 data_array.data0\[1\]\[41\] VGND VGND VPWR VPWR net1965 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold325 data_array.data1\[0\]\[24\] VGND VGND VPWR VPWR net1976 sky130_fd_sc_hd__dlygate4sd3_1
Xhold336 data_array.data0\[4\]\[41\] VGND VGND VPWR VPWR net1987 sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 data_array.data0\[0\]\[62\] VGND VGND VPWR VPWR net1998 sky130_fd_sc_hd__dlygate4sd3_1
Xhold358 data_array.data1\[0\]\[45\] VGND VGND VPWR VPWR net2009 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09931_ net1105 net3620 net370 VGND VGND VPWR VPWR _01680_ sky130_fd_sc_hd__mux2_1
Xhold369 data_array.data0\[4\]\[63\] VGND VGND VPWR VPWR net2020 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout805 net806 VGND VGND VPWR VPWR net805 sky130_fd_sc_hd__clkbuf_8
Xfanout816 _05359_ VGND VGND VPWR VPWR net816 sky130_fd_sc_hd__clkbuf_4
X_09862_ net1020 net2596 net379 VGND VGND VPWR VPWR _01612_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_74_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout838 net844 VGND VGND VPWR VPWR net838 sky130_fd_sc_hd__buf_8
Xfanout849 net853 VGND VGND VPWR VPWR net849 sky130_fd_sc_hd__buf_4
XFILLER_100_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1003 data_array.data1\[9\]\[62\] VGND VGND VPWR VPWR net2654 sky130_fd_sc_hd__dlygate4sd3_1
X_08813_ net1918 net993 net447 VGND VGND VPWR VPWR _00571_ sky130_fd_sc_hd__mux2_1
Xhold1014 data_array.data1\[5\]\[44\] VGND VGND VPWR VPWR net2665 sky130_fd_sc_hd__dlygate4sd3_1
X_09793_ net1036 net3262 net387 VGND VGND VPWR VPWR _01544_ sky130_fd_sc_hd__mux2_1
Xhold1025 tag_array.tag1\[8\]\[23\] VGND VGND VPWR VPWR net2676 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1036 data_array.data0\[6\]\[5\] VGND VGND VPWR VPWR net2687 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1047 tag_array.tag1\[12\]\[19\] VGND VGND VPWR VPWR net2698 sky130_fd_sc_hd__dlygate4sd3_1
X_05956_ net134 net1151 _03430_ _03431_ VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__a22o_1
X_08744_ net747 net3603 net460 VGND VGND VPWR VPWR _00503_ sky130_fd_sc_hd__mux2_1
Xhold1058 tag_array.tag0\[10\]\[10\] VGND VGND VPWR VPWR net2709 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1069 data_array.data1\[14\]\[15\] VGND VGND VPWR VPWR net2720 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08675_ net724 net3551 net500 VGND VGND VPWR VPWR _00434_ sky130_fd_sc_hd__mux2_1
X_05887_ net108 net1154 _03384_ _03385_ VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__a22o_1
XFILLER_81_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07626_ net1170 _04845_ _04849_ net1218 VGND VGND VPWR VPWR _04851_ sky130_fd_sc_hd__a22o_1
XFILLER_53_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07557_ data_array.data1\[1\]\[10\] net1606 net1510 data_array.data1\[2\]\[10\] VGND
+ VGND VPWR VPWR _04788_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_33_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_33_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_157_3373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06508_ tag_array.tag1\[1\]\[4\] net1552 net1456 tag_array.tag1\[2\]\[4\] VGND VGND
+ VPWR VPWR _03834_ sky130_fd_sc_hd__a22o_1
XFILLER_22_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_3384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07488_ data_array.data1\[4\]\[4\] net1393 net1299 data_array.data1\[7\]\[4\] _04724_
+ VGND VGND VPWR VPWR _04725_ sky130_fd_sc_hd__a221o_1
XFILLER_21_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06439_ _03770_ _03771_ VGND VGND VPWR VPWR _00145_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_118_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09227_ net770 net2937 net647 VGND VGND VPWR VPWR _00981_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_118_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09158_ net908 net4201 net567 VGND VGND VPWR VPWR _00912_ sky130_fd_sc_hd__mux2_1
XFILLER_5_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08109_ net1635 _05283_ _05287_ net1209 VGND VGND VPWR VPWR _05290_ sky130_fd_sc_hd__a22o_1
XFILLER_108_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09089_ net928 net3815 net411 VGND VGND VPWR VPWR _00843_ sky130_fd_sc_hd__mux2_1
X_11120_ net1039 net4067 net543 VGND VGND VPWR VPWR _02863_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_131_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold870 data_array.data0\[12\]\[45\] VGND VGND VPWR VPWR net2521 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_131_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold881 data_array.data0\[1\]\[38\] VGND VGND VPWR VPWR net2532 sky130_fd_sc_hd__dlygate4sd3_1
X_11051_ net1738 net1058 net330 VGND VGND VPWR VPWR _02794_ sky130_fd_sc_hd__mux2_1
XFILLER_104_952 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold892 data_array.data0\[5\]\[24\] VGND VGND VPWR VPWR net2543 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_567 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10002_ net1079 net3243 net556 VGND VGND VPWR VPWR _01751_ sky130_fd_sc_hd__mux2_1
XFILLER_27_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2260 data_array.data1\[10\]\[8\] VGND VGND VPWR VPWR net3911 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2271 data_array.data1\[12\]\[12\] VGND VGND VPWR VPWR net3922 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2282 data_array.data1\[11\]\[18\] VGND VGND VPWR VPWR net3933 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2293 tag_array.tag1\[6\]\[5\] VGND VGND VPWR VPWR net3944 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1570 data_array.data1\[5\]\[31\] VGND VGND VPWR VPWR net3221 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1581 data_array.data0\[2\]\[41\] VGND VGND VPWR VPWR net3232 sky130_fd_sc_hd__dlygate4sd3_1
X_11953_ clknet_leaf_229_clk _00761_ VGND VGND VPWR VPWR data_array.data0\[4\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1592 data_array.data1\[13\]\[8\] VGND VGND VPWR VPWR net3243 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_28_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10904_ net870 net3511 net523 VGND VGND VPWR VPWR _02649_ sky130_fd_sc_hd__mux2_1
XFILLER_83_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11884_ clknet_leaf_9_clk _00692_ VGND VGND VPWR VPWR data_array.data0\[5\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_13623_ clknet_leaf_90_clk _02252_ VGND VGND VPWR VPWR data_array.data0\[9\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
X_10835_ net2645 net890 net503 VGND VGND VPWR VPWR _02580_ sky130_fd_sc_hd__mux2_1
XFILLER_13_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_24_clk clknet_5_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_8
X_13554_ clknet_leaf_4_clk _02183_ VGND VGND VPWR VPWR data_array.data1\[0\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10766_ net908 net4290 net491 VGND VGND VPWR VPWR _02511_ sky130_fd_sc_hd__mux2_1
XFILLER_160_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12505_ clknet_leaf_238_clk _01199_ VGND VGND VPWR VPWR data_array.data1\[9\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
X_10697_ net2083 net930 net479 VGND VGND VPWR VPWR _02442_ sky130_fd_sc_hd__mux2_1
X_13485_ clknet_leaf_144_clk _02115_ VGND VGND VPWR VPWR tag_array.tag0\[15\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_157_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12436_ clknet_leaf_220_clk _01130_ VGND VGND VPWR VPWR data_array.data0\[14\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12367_ clknet_leaf_62_clk _00043_ VGND VGND VPWR VPWR data_array.rdata0\[49\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_39_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14106_ clknet_leaf_15_clk _02735_ VGND VGND VPWR VPWR data_array.data0\[1\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11318_ net1021 net2955 net796 VGND VGND VPWR VPWR _03061_ sky130_fd_sc_hd__mux2_1
X_12298_ clknet_leaf_136_clk _01056_ VGND VGND VPWR VPWR tag_array.tag1\[12\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_56_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11249_ net1035 net3541 net681 VGND VGND VPWR VPWR _02992_ sky130_fd_sc_hd__mux2_1
X_14037_ clknet_leaf_201_clk _02666_ VGND VGND VPWR VPWR data_array.data1\[6\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_79_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_52_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05810_ _03156_ _03158_ _03203_ _03214_ VGND VGND VPWR VPWR _03327_ sky130_fd_sc_hd__or4_1
X_06790_ net1178 _04085_ _04089_ net1226 VGND VGND VPWR VPWR _04091_ sky130_fd_sc_hd__a22o_1
X_05741_ fsm.tag_out1\[1\] net31 VGND VGND VPWR VPWR _03258_ sky130_fd_sc_hd__and2b_1
XFILLER_48_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08460_ net157 net92 net1648 VGND VGND VPWR VPWR _05543_ sky130_fd_sc_hd__mux2_1
X_05672_ fsm.tag_out0\[15\] net15 VGND VGND VPWR VPWR _03189_ sky130_fd_sc_hd__and2b_1
X_07411_ data_array.data0\[0\]\[61\] net1357 net1263 data_array.data0\[3\]\[61\] _04654_
+ VGND VGND VPWR VPWR _04655_ sky130_fd_sc_hd__a221o_1
XFILLER_23_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08391_ net131 net66 net1639 VGND VGND VPWR VPWR _05497_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_15_clk clknet_5_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_8
X_07342_ data_array.data0\[13\]\[55\] net1534 net1438 data_array.data0\[14\]\[55\]
+ VGND VGND VPWR VPWR _04592_ sky130_fd_sc_hd__a22o_1
XFILLER_177_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07273_ net1630 _04523_ _04527_ net1204 VGND VGND VPWR VPWR _04530_ sky130_fd_sc_hd__a22o_1
X_09012_ net2435 net976 net422 VGND VGND VPWR VPWR _00767_ sky130_fd_sc_hd__mux2_1
X_06224_ tag_array.tag0\[9\]\[3\] net1564 net1468 tag_array.tag0\[10\]\[3\] VGND VGND
+ VPWR VPWR _03576_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_152_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold100 data_array.data0\[2\]\[2\] VGND VGND VPWR VPWR net1751 sky130_fd_sc_hd__dlygate4sd3_1
X_06155_ tag_array.valid0\[9\] net1597 net1501 tag_array.valid0\[10\] VGND VGND VPWR
+ VPWR _03512_ sky130_fd_sc_hd__a22o_1
Xhold111 data_array.data1\[1\]\[26\] VGND VGND VPWR VPWR net1762 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold122 data_array.data0\[2\]\[10\] VGND VGND VPWR VPWR net1773 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold133 tag_array.tag1\[1\]\[1\] VGND VGND VPWR VPWR net1784 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold144 tag_array.tag1\[4\]\[10\] VGND VGND VPWR VPWR net1795 sky130_fd_sc_hd__dlygate4sd3_1
X_06086_ data_array.rdata0\[1\] net1134 net1112 data_array.rdata1\[1\] VGND VGND VPWR
+ VPWR net274 sky130_fd_sc_hd__a22o_1
Xhold155 data_array.data0\[4\]\[31\] VGND VGND VPWR VPWR net1806 sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 tag_array.tag1\[4\]\[19\] VGND VGND VPWR VPWR net1817 sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 data_array.data1\[4\]\[56\] VGND VGND VPWR VPWR net1828 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold188 data_array.data0\[4\]\[51\] VGND VGND VPWR VPWR net1839 sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 data_array.data0\[1\]\[15\] VGND VGND VPWR VPWR net1850 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout602 net604 VGND VGND VPWR VPWR net602 sky130_fd_sc_hd__buf_4
X_09914_ net752 net3462 net603 VGND VGND VPWR VPWR _01664_ sky130_fd_sc_hd__mux2_1
Xfanout613 net614 VGND VGND VPWR VPWR net613 sky130_fd_sc_hd__buf_4
Xfanout624 _05565_ VGND VGND VPWR VPWR net624 sky130_fd_sc_hd__buf_4
Xfanout635 net636 VGND VGND VPWR VPWR net635 sky130_fd_sc_hd__buf_4
XFILLER_99_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout646 net647 VGND VGND VPWR VPWR net646 sky130_fd_sc_hd__buf_4
Xfanout657 net660 VGND VGND VPWR VPWR net657 sky130_fd_sc_hd__buf_2
X_09845_ net1088 net2454 net380 VGND VGND VPWR VPWR _01595_ sky130_fd_sc_hd__mux2_1
XFILLER_58_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout668 net670 VGND VGND VPWR VPWR net668 sky130_fd_sc_hd__buf_4
Xfanout679 _05548_ VGND VGND VPWR VPWR net679 sky130_fd_sc_hd__clkbuf_4
XFILLER_85_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09776_ net1106 net4029 net386 VGND VGND VPWR VPWR _01527_ sky130_fd_sc_hd__mux2_1
X_06988_ net1216 _04265_ _04269_ net1168 VGND VGND VPWR VPWR _04271_ sky130_fd_sc_hd__a22o_1
XFILLER_37_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08727_ net1808 net714 net476 VGND VGND VPWR VPWR _00486_ sky130_fd_sc_hd__mux2_1
X_05939_ data_array.rdata0\[36\] net1659 net1149 VGND VGND VPWR VPWR _03420_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_159_3413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_159_3424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ net791 net2853 net496 VGND VGND VPWR VPWR _00417_ sky130_fd_sc_hd__mux2_1
XFILLER_41_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07609_ data_array.data1\[4\]\[15\] net1394 net1300 data_array.data1\[7\]\[15\] _04834_
+ VGND VGND VPWR VPWR _04835_ sky130_fd_sc_hd__a221o_1
X_08589_ _05377_ net3592 net530 VGND VGND VPWR VPWR _00348_ sky130_fd_sc_hd__mux2_1
X_10620_ net2054 net980 net466 VGND VGND VPWR VPWR _02365_ sky130_fd_sc_hd__mux2_1
XFILLER_169_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10551_ net1001 net3971 net454 VGND VGND VPWR VPWR _02296_ sky130_fd_sc_hd__mux2_1
XFILLER_139_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10482_ net1019 net4372 net347 VGND VGND VPWR VPWR _02227_ sky130_fd_sc_hd__mux2_1
X_13270_ clknet_leaf_46_clk _01900_ VGND VGND VPWR VPWR data_array.data0\[11\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_133_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12221_ clknet_leaf_183_clk _00174_ VGND VGND VPWR VPWR fsm.tag_out1\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12152_ clknet_leaf_158_clk _00960_ VGND VGND VPWR VPWR tag_array.tag0\[13\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11103_ net1107 net3275 net541 VGND VGND VPWR VPWR _02846_ sky130_fd_sc_hd__mux2_1
X_12083_ clknet_leaf_39_clk _00891_ VGND VGND VPWR VPWR data_array.data1\[14\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_150_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_771 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11034_ net2133 net866 net338 VGND VGND VPWR VPWR _02778_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_34_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2090 data_array.data0\[5\]\[37\] VGND VGND VPWR VPWR net3741 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12985_ clknet_leaf_230_clk _01679_ VGND VGND VPWR VPWR data_array.data0\[3\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_11936_ clknet_leaf_111_clk _00744_ VGND VGND VPWR VPWR data_array.data0\[4\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11867_ clknet_leaf_210_clk _00675_ VGND VGND VPWR VPWR data_array.data0\[5\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_13606_ clknet_leaf_38_clk _02235_ VGND VGND VPWR VPWR data_array.data0\[9\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_10818_ net3114 net958 net509 VGND VGND VPWR VPWR _02563_ sky130_fd_sc_hd__mux2_1
XFILLER_159_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11798_ clknet_leaf_230_clk _00606_ VGND VGND VPWR VPWR data_array.data0\[7\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_13537_ clknet_leaf_7_clk _02166_ VGND VGND VPWR VPWR data_array.data1\[0\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
X_10749_ net978 net4612 net497 VGND VGND VPWR VPWR _02494_ sky130_fd_sc_hd__mux2_1
XFILLER_174_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13468_ clknet_leaf_190_clk _02098_ VGND VGND VPWR VPWR tag_array.tag0\[1\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_127_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12419_ clknet_leaf_219_clk _01113_ VGND VGND VPWR VPWR data_array.data0\[14\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_93_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13399_ clknet_leaf_67_clk _02029_ VGND VGND VPWR VPWR data_array.data1\[8\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput205 net205 VGND VGND VPWR VPWR cpu_rdata[46] sky130_fd_sc_hd__buf_4
XFILLER_142_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput216 net216 VGND VGND VPWR VPWR cpu_rdata[56] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_93_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput227 net227 VGND VGND VPWR VPWR cpu_rdata[8] sky130_fd_sc_hd__buf_2
XFILLER_142_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput238 net238 VGND VGND VPWR VPWR mem_addr[17] sky130_fd_sc_hd__buf_2
Xoutput249 net249 VGND VGND VPWR VPWR mem_addr[27] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_34_Left_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07960_ data_array.data1\[5\]\[47\] net1588 net1492 data_array.data1\[6\]\[47\] VGND
+ VGND VPWR VPWR _05154_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_4_clk clknet_5_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_71_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06911_ net1180 _04195_ _04199_ net1228 VGND VGND VPWR VPWR _04201_ sky130_fd_sc_hd__a22o_1
XFILLER_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07891_ _05090_ _05091_ VGND VGND VPWR VPWR _00098_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_155_Right_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09630_ net769 net4192 net615 VGND VGND VPWR VPWR _01382_ sky130_fd_sc_hd__mux2_1
X_06842_ data_array.data0\[1\]\[9\] net1580 net1484 data_array.data0\[2\]\[9\] VGND
+ VGND VPWR VPWR _04138_ sky130_fd_sc_hd__a22o_1
X_09561_ net1106 net4577 net394 VGND VGND VPWR VPWR _01313_ sky130_fd_sc_hd__mux2_1
X_06773_ data_array.data0\[4\]\[3\] net1377 net1283 data_array.data0\[7\]\[3\] _04074_
+ VGND VGND VPWR VPWR _04075_ sky130_fd_sc_hd__a221o_1
X_08512_ net821 net811 net854 _05577_ VGND VGND VPWR VPWR _05579_ sky130_fd_sc_hd__or4b_1
XFILLER_82_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05724_ _03237_ _03238_ _03239_ _03240_ VGND VGND VPWR VPWR _03241_ sky130_fd_sc_hd__or4_1
XFILLER_36_563 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09492_ net761 net3619 net626 VGND VGND VPWR VPWR _01245_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_43_Left_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08443_ net1124 _05531_ VGND VGND VPWR VPWR _05532_ sky130_fd_sc_hd__and2_1
X_05655_ fsm.tag_out0\[21\] net21 VGND VGND VPWR VPWR _03172_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_137_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08374_ net1127 _05485_ VGND VGND VPWR VPWR _05486_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_154_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07325_ data_array.data0\[12\]\[53\] net1332 net1238 data_array.data0\[15\]\[53\]
+ _04576_ VGND VGND VPWR VPWR _04577_ sky130_fd_sc_hd__a221o_1
XFILLER_139_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_5_18__f_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_5_18__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_17_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07256_ data_array.data0\[5\]\[47\] net1578 net1482 data_array.data0\[6\]\[47\] VGND
+ VGND VPWR VPWR _04514_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_30_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06207_ net1181 _03555_ _03559_ net1229 VGND VGND VPWR VPWR _03561_ sky130_fd_sc_hd__a22o_1
XFILLER_180_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07187_ _04450_ _04451_ VGND VGND VPWR VPWR _00034_ sky130_fd_sc_hd__or2_1
XFILLER_155_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_52_Left_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06138_ data_array.rdata0\[53\] net1134 net1112 data_array.rdata1\[53\] VGND VGND
+ VPWR VPWR net311 sky130_fd_sc_hd__a22o_1
XFILLER_132_332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06069_ net1163 net17 fsm.tag_out1\[17\] net1133 VGND VGND VPWR VPWR _03498_ sky130_fd_sc_hd__a22o_1
XFILLER_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout410 net417 VGND VGND VPWR VPWR net410 sky130_fd_sc_hd__clkbuf_8
Xfanout1408 net1422 VGND VGND VPWR VPWR net1408 sky130_fd_sc_hd__clkbuf_2
XFILLER_160_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1419 net1420 VGND VGND VPWR VPWR net1419 sky130_fd_sc_hd__clkbuf_4
Xfanout421 net425 VGND VGND VPWR VPWR net421 sky130_fd_sc_hd__buf_4
Xfanout432 net433 VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__buf_4
Xfanout443 net449 VGND VGND VPWR VPWR net443 sky130_fd_sc_hd__clkbuf_8
Xfanout454 net459 VGND VGND VPWR VPWR net454 sky130_fd_sc_hd__clkbuf_4
XFILLER_87_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout465 _05604_ VGND VGND VPWR VPWR net465 sky130_fd_sc_hd__clkbuf_4
Xfanout476 net477 VGND VGND VPWR VPWR net476 sky130_fd_sc_hd__buf_4
Xfanout487 net488 VGND VGND VPWR VPWR net487 sky130_fd_sc_hd__buf_4
X_09828_ net897 net2842 net386 VGND VGND VPWR VPWR _01579_ sky130_fd_sc_hd__mux2_1
XFILLER_59_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_122_Right_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout498 net499 VGND VGND VPWR VPWR net498 sky130_fd_sc_hd__buf_2
XFILLER_171_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09759_ net2868 net750 net672 VGND VGND VPWR VPWR _01511_ sky130_fd_sc_hd__mux2_1
XFILLER_39_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_126_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_61_Left_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ clknet_leaf_144_clk _01464_ VGND VGND VPWR VPWR tag_array.tag0\[6\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_161_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_174_3708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ clknet_leaf_153_clk _00529_ VGND VGND VPWR VPWR tag_array.tag0\[9\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_14440_ clknet_leaf_91_clk _03063_ VGND VGND VPWR VPWR data_array.data1\[7\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11652_ clknet_leaf_186_clk _00460_ VGND VGND VPWR VPWR tag_array.tag1\[2\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10603_ net1725 net1051 net472 VGND VGND VPWR VPWR _02348_ sky130_fd_sc_hd__mux2_1
X_14371_ clknet_leaf_221_clk _02994_ VGND VGND VPWR VPWR data_array.data1\[10\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_11583_ clknet_leaf_189_clk _00391_ VGND VGND VPWR VPWR tag_array.tag1\[5\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13322_ clknet_leaf_38_clk _01952_ VGND VGND VPWR VPWR data_array.data0\[10\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_10534_ net1070 net3458 net463 VGND VGND VPWR VPWR _02279_ sky130_fd_sc_hd__mux2_1
XFILLER_7_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_70_Left_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10465_ net1084 net2840 net344 VGND VGND VPWR VPWR _02210_ sky130_fd_sc_hd__mux2_1
X_13253_ clknet_leaf_240_clk _01883_ VGND VGND VPWR VPWR data_array.data0\[11\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12204_ clknet_leaf_151_clk _00133_ VGND VGND VPWR VPWR fsm.tag_out0\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_136_682 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10396_ net1741 net1070 net671 VGND VGND VPWR VPWR _02142_ sky130_fd_sc_hd__mux2_1
X_13184_ clknet_leaf_215_clk _00077_ VGND VGND VPWR VPWR data_array.rdata1\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12135_ clknet_leaf_159_clk _00943_ VGND VGND VPWR VPWR tag_array.tag0\[12\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_111_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12066_ clknet_leaf_85_clk _00874_ VGND VGND VPWR VPWR data_array.data1\[14\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11017_ net2113 net932 _03132_ VGND VGND VPWR VPWR _02761_ sky130_fd_sc_hd__mux2_1
XFILLER_38_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12968_ clknet_leaf_144_clk _01662_ VGND VGND VPWR VPWR tag_array.tag0\[4\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11919_ clknet_leaf_237_clk _00727_ VGND VGND VPWR VPWR data_array.data0\[5\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
X_12899_ clknet_leaf_46_clk _01593_ VGND VGND VPWR VPWR data_array.data0\[13\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_178_549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_109_Left_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07110_ _04380_ _04381_ VGND VGND VPWR VPWR _00026_ sky130_fd_sc_hd__or2_1
X_08090_ data_array.data1\[9\]\[59\] net1572 net1476 data_array.data1\[10\]\[59\]
+ VGND VGND VPWR VPWR _05272_ sky130_fd_sc_hd__a22o_1
XFILLER_174_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload20 clknet_leaf_270_clk VGND VGND VPWR VPWR clkload20/Y sky130_fd_sc_hd__inv_8
X_07041_ data_array.data0\[4\]\[27\] net1365 net1271 data_array.data0\[7\]\[27\] _04318_
+ VGND VGND VPWR VPWR _04319_ sky130_fd_sc_hd__a221o_1
Xclkload31 clknet_leaf_11_clk VGND VGND VPWR VPWR clkload31/Y sky130_fd_sc_hd__clkinv_2
Xclkload42 clknet_leaf_22_clk VGND VGND VPWR VPWR clkload42/Y sky130_fd_sc_hd__bufinv_16
Xclkload53 clknet_leaf_251_clk VGND VGND VPWR VPWR clkload53/X sky130_fd_sc_hd__clkbuf_4
Xclkload64 clknet_leaf_242_clk VGND VGND VPWR VPWR clkload64/Y sky130_fd_sc_hd__clkinv_4
XFILLER_173_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload75 clknet_leaf_47_clk VGND VGND VPWR VPWR clkload75/Y sky130_fd_sc_hd__bufinv_16
Xclkload86 clknet_leaf_46_clk VGND VGND VPWR VPWR clkload86/Y sky130_fd_sc_hd__clkinv_2
Xclkload97 clknet_leaf_59_clk VGND VGND VPWR VPWR clkload97/Y sky130_fd_sc_hd__inv_8
XFILLER_173_1034 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08992_ net2593 net1058 net420 VGND VGND VPWR VPWR _00747_ sky130_fd_sc_hd__mux2_1
Xhold2804 tag_array.tag0\[1\]\[1\] VGND VGND VPWR VPWR net4455 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2815 data_array.data0\[15\]\[22\] VGND VGND VPWR VPWR net4466 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_141_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2826 data_array.data1\[6\]\[45\] VGND VGND VPWR VPWR net4477 sky130_fd_sc_hd__dlygate4sd3_1
X_07943_ data_array.data1\[4\]\[45\] net1350 net1256 data_array.data1\[7\]\[45\] _05138_
+ VGND VGND VPWR VPWR _05139_ sky130_fd_sc_hd__a221o_1
Xhold2837 data_array.data0\[6\]\[29\] VGND VGND VPWR VPWR net4488 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2848 data_array.data0\[9\]\[28\] VGND VGND VPWR VPWR net4499 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_147_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2859 data_array.data0\[3\]\[11\] VGND VGND VPWR VPWR net4510 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_68_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07874_ data_array.data1\[13\]\[39\] net1538 net1442 data_array.data1\[14\]\[39\]
+ VGND VGND VPWR VPWR _05076_ sky130_fd_sc_hd__a22o_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09613_ net897 net2755 net394 VGND VGND VPWR VPWR _01365_ sky130_fd_sc_hd__mux2_1
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06825_ data_array.data0\[13\]\[8\] net1536 net1440 data_array.data0\[14\]\[8\] VGND
+ VGND VPWR VPWR _04122_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_108_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09544_ net751 net3309 net619 VGND VGND VPWR VPWR _01297_ sky130_fd_sc_hd__mux2_1
X_06756_ net1188 _04053_ _04057_ net1614 VGND VGND VPWR VPWR _04060_ sky130_fd_sc_hd__a22o_1
XFILLER_37_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05707_ net32 fsm.tag_out0\[2\] VGND VGND VPWR VPWR _03224_ sky130_fd_sc_hd__and2b_1
X_09475_ net729 net3599 net658 VGND VGND VPWR VPWR _01228_ sky130_fd_sc_hd__mux2_1
XFILLER_34_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06687_ tag_array.tag1\[12\]\[20\] net1368 net1274 tag_array.tag1\[15\]\[20\] _03996_
+ VGND VGND VPWR VPWR _03997_ sky130_fd_sc_hd__a221o_1
XFILLER_180_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08426_ net2273 net909 net687 VGND VGND VPWR VPWR _00271_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_121_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05638_ net11 fsm.tag_out0\[12\] VGND VGND VPWR VPWR _03155_ sky130_fd_sc_hd__xor2_1
XFILLER_180_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08357_ net2064 net1002 net689 VGND VGND VPWR VPWR _00248_ sky130_fd_sc_hd__mux2_1
XFILLER_133_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload3 clknet_5_6__leaf_clk VGND VGND VPWR VPWR clkload3/X sky130_fd_sc_hd__clkbuf_8
X_07308_ _04560_ _04561_ VGND VGND VPWR VPWR _00046_ sky130_fd_sc_hd__or2_1
XFILLER_138_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08288_ net2056 net1092 net691 VGND VGND VPWR VPWR _00225_ sky130_fd_sc_hd__mux2_1
XFILLER_165_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07239_ data_array.data0\[4\]\[45\] net1344 net1250 data_array.data0\[7\]\[45\] _04498_
+ VGND VGND VPWR VPWR _04499_ sky130_fd_sc_hd__a221o_1
X_10250_ net745 net2397 net595 VGND VGND VPWR VPWR _01997_ sky130_fd_sc_hd__mux2_1
X_10181_ net1081 net3823 net360 VGND VGND VPWR VPWR _01928_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_167_3567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_167_3578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1205 net1206 VGND VGND VPWR VPWR net1205 sky130_fd_sc_hd__buf_4
XFILLER_59_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1216 net1217 VGND VGND VPWR VPWR net1216 sky130_fd_sc_hd__buf_4
XFILLER_132_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1227 net1228 VGND VGND VPWR VPWR net1227 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_184_3892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1238 net1240 VGND VGND VPWR VPWR net1238 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_128_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1249 net1251 VGND VGND VPWR VPWR net1249 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_128_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13940_ clknet_leaf_78_clk _02569_ VGND VGND VPWR VPWR data_array.data1\[4\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13871_ clknet_leaf_240_clk _02500_ VGND VGND VPWR VPWR data_array.data1\[3\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12822_ clknet_leaf_98_clk _01516_ VGND VGND VPWR VPWR tag_array.tag1\[0\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12753_ clknet_leaf_158_clk _01447_ VGND VGND VPWR VPWR tag_array.tag0\[5\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11704_ clknet_leaf_232_clk _00512_ VGND VGND VPWR VPWR tag_array.tag1\[15\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_91_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12684_ clknet_leaf_170_clk _01378_ VGND VGND VPWR VPWR tag_array.tag0\[8\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_14423_ clknet_leaf_82_clk _03046_ VGND VGND VPWR VPWR data_array.data1\[7\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_11635_ clknet_leaf_99_clk _00443_ VGND VGND VPWR VPWR tag_array.tag1\[2\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14354_ clknet_leaf_68_clk _02977_ VGND VGND VPWR VPWR data_array.data1\[10\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_11566_ clknet_leaf_132_clk _00374_ VGND VGND VPWR VPWR tag_array.tag1\[5\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13305_ clknet_leaf_50_clk _01935_ VGND VGND VPWR VPWR data_array.data0\[10\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_156_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10517_ net876 net4501 net346 VGND VGND VPWR VPWR _02262_ sky130_fd_sc_hd__mux2_1
X_14285_ clknet_leaf_199_clk _02914_ VGND VGND VPWR VPWR data_array.data1\[11\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11497_ clknet_leaf_172_clk _00305_ VGND VGND VPWR VPWR tag_array.valid1\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_90_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13236_ clknet_leaf_60_clk _01866_ VGND VGND VPWR VPWR data_array.data0\[11\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_10448_ net2038 net862 net671 VGND VGND VPWR VPWR _02194_ sky130_fd_sc_hd__mux2_1
XFILLER_171_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13167_ clknet_leaf_68_clk _00108_ VGND VGND VPWR VPWR data_array.rdata1\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_69_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10379_ net353 net2635 net569 VGND VGND VPWR VPWR _02125_ sky130_fd_sc_hd__mux2_1
XFILLER_111_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12118_ clknet_leaf_159_clk _00926_ VGND VGND VPWR VPWR tag_array.tag0\[12\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_85_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13098_ clknet_leaf_56_clk _01792_ VGND VGND VPWR VPWR data_array.data1\[13\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
X_12049_ clknet_leaf_52_clk _00857_ VGND VGND VPWR VPWR data_array.data0\[6\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_65_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_88_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06610_ tag_array.tag1\[8\]\[13\] net1420 net1326 tag_array.tag1\[11\]\[13\] _03926_
+ VGND VGND VPWR VPWR _03927_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_49_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07590_ data_array.data1\[5\]\[13\] net1550 net1454 data_array.data1\[6\]\[13\] VGND
+ VGND VPWR VPWR _04818_ sky130_fd_sc_hd__a22o_1
XFILLER_80_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06541_ tag_array.tag1\[5\]\[7\] net1610 net1514 tag_array.tag1\[6\]\[7\] VGND VGND
+ VPWR VPWR _03864_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_66_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09260_ net741 net2415 net577 VGND VGND VPWR VPWR _01014_ sky130_fd_sc_hd__mux2_1
X_06472_ _03800_ _03801_ VGND VGND VPWR VPWR _00156_ sky130_fd_sc_hd__or2_2
XFILLER_179_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_117_Left_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08211_ net773 net2347 net804 VGND VGND VPWR VPWR _00201_ sky130_fd_sc_hd__mux2_1
X_09191_ net716 net2975 net628 VGND VGND VPWR VPWR _00945_ sky130_fd_sc_hd__mux2_1
XFILLER_159_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08142_ net1196 _05313_ _05317_ net1623 VGND VGND VPWR VPWR _05320_ sky130_fd_sc_hd__a22o_1
XFILLER_140_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload120 clknet_leaf_76_clk VGND VGND VPWR VPWR clkload120/Y sky130_fd_sc_hd__clkinv_8
X_08073_ data_array.data1\[8\]\[57\] net1347 net1253 data_array.data1\[11\]\[57\]
+ _05256_ VGND VGND VPWR VPWR _05257_ sky130_fd_sc_hd__a221o_1
Xclkload131 clknet_leaf_87_clk VGND VGND VPWR VPWR clkload131/X sky130_fd_sc_hd__clkbuf_4
XFILLER_146_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload142 clknet_leaf_207_clk VGND VGND VPWR VPWR clkload142/X sky130_fd_sc_hd__clkbuf_8
X_07024_ data_array.data0\[8\]\[26\] net1338 net1244 data_array.data0\[11\]\[26\]
+ _04302_ VGND VGND VPWR VPWR _04303_ sky130_fd_sc_hd__a221o_1
Xclkload153 clknet_leaf_230_clk VGND VGND VPWR VPWR clkload153/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload164 clknet_leaf_202_clk VGND VGND VPWR VPWR clkload164/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload175 clknet_leaf_200_clk VGND VGND VPWR VPWR clkload175/Y sky130_fd_sc_hd__clkinv_2
Xclkload186 clknet_leaf_187_clk VGND VGND VPWR VPWR clkload186/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_149_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload197 clknet_leaf_106_clk VGND VGND VPWR VPWR clkload197/Y sky130_fd_sc_hd__bufinv_16
XFILLER_88_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_126_Left_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2601 data_array.data0\[13\]\[45\] VGND VGND VPWR VPWR net4252 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_142_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2612 data_array.data1\[5\]\[14\] VGND VGND VPWR VPWR net4263 sky130_fd_sc_hd__dlygate4sd3_1
X_08975_ net866 net4321 net429 VGND VGND VPWR VPWR _00731_ sky130_fd_sc_hd__mux2_1
Xhold2623 data_array.data0\[11\]\[31\] VGND VGND VPWR VPWR net4274 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2634 data_array.data0\[11\]\[29\] VGND VGND VPWR VPWR net4285 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1900 tag_array.tag1\[3\]\[17\] VGND VGND VPWR VPWR net3551 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2645 data_array.data1\[11\]\[32\] VGND VGND VPWR VPWR net4296 sky130_fd_sc_hd__dlygate4sd3_1
X_07926_ data_array.data1\[8\]\[44\] net1398 net1304 data_array.data1\[11\]\[44\]
+ _05122_ VGND VGND VPWR VPWR _05123_ sky130_fd_sc_hd__a221o_1
Xhold2656 tag_array.tag1\[7\]\[2\] VGND VGND VPWR VPWR net4307 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1911 tag_array.tag0\[3\]\[17\] VGND VGND VPWR VPWR net3562 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2667 data_array.data0\[6\]\[41\] VGND VGND VPWR VPWR net4318 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 tag_array.valid1\[10\] VGND VGND VPWR VPWR net1699 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1922 tag_array.tag0\[1\]\[15\] VGND VGND VPWR VPWR net3573 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1933 tag_array.tag1\[7\]\[20\] VGND VGND VPWR VPWR net3584 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 tag_array.valid0\[5\] VGND VGND VPWR VPWR net1710 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2678 data_array.data0\[10\]\[29\] VGND VGND VPWR VPWR net4329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2689 data_array.data1\[5\]\[40\] VGND VGND VPWR VPWR net4340 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_162_3475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1944 data_array.data1\[3\]\[56\] VGND VGND VPWR VPWR net3595 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1955 data_array.data0\[10\]\[60\] VGND VGND VPWR VPWR net3606 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_21_1029 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07857_ net1218 _05055_ _05059_ net1170 VGND VGND VPWR VPWR _05061_ sky130_fd_sc_hd__a22o_1
XFILLER_56_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1966 data_array.data1\[15\]\[22\] VGND VGND VPWR VPWR net3617 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1977 data_array.data1\[6\]\[44\] VGND VGND VPWR VPWR net3628 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1988 data_array.data1\[10\]\[35\] VGND VGND VPWR VPWR net3639 sky130_fd_sc_hd__dlygate4sd3_1
X_06808_ data_array.data0\[12\]\[6\] net1331 net1237 data_array.data0\[15\]\[6\] _04106_
+ VGND VGND VPWR VPWR _04107_ sky130_fd_sc_hd__a221o_1
XFILLER_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_123_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1999 data_array.data0\[3\]\[9\] VGND VGND VPWR VPWR net3650 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_71_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07788_ data_array.data1\[1\]\[31\] net1572 net1476 data_array.data1\[2\]\[31\] VGND
+ VGND VPWR VPWR _04998_ sky130_fd_sc_hd__a22o_1
X_09527_ net719 net2993 net621 VGND VGND VPWR VPWR _01280_ sky130_fd_sc_hd__mux2_1
XFILLER_24_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06739_ data_array.data0\[1\]\[0\] net1555 net1459 data_array.data0\[2\]\[0\] VGND
+ VGND VPWR VPWR _04044_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_135_Left_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09458_ net819 net3762 _05564_ VGND VGND VPWR VPWR _01211_ sky130_fd_sc_hd__mux2_1
X_08409_ net138 net73 net1639 VGND VGND VPWR VPWR _05509_ sky130_fd_sc_hd__mux2_1
X_09389_ net1110 net2836 net584 VGND VGND VPWR VPWR _01142_ sky130_fd_sc_hd__mux2_1
X_11420_ clknet_leaf_61_clk _00230_ VGND VGND VPWR VPWR data_array.data0\[0\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_530 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11351_ net890 net3751 net796 VGND VGND VPWR VPWR _03094_ sky130_fd_sc_hd__mux2_1
XFILLER_125_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_169_3607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_169_3618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10302_ net2245 net952 net634 VGND VGND VPWR VPWR _02049_ sky130_fd_sc_hd__mux2_1
XFILLER_152_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14070_ clknet_leaf_261_clk _02699_ VGND VGND VPWR VPWR data_array.data1\[6\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
X_11282_ net900 net3284 net677 VGND VGND VPWR VPWR _03025_ sky130_fd_sc_hd__mux2_1
X_13021_ clknet_leaf_114_clk _01715_ VGND VGND VPWR VPWR data_array.data0\[3\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10233_ net873 net3883 net358 VGND VGND VPWR VPWR _01980_ sky130_fd_sc_hd__mux2_1
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1002 net1003 VGND VGND VPWR VPWR net1002 sky130_fd_sc_hd__clkbuf_2
X_10164_ net889 net4515 net363 VGND VGND VPWR VPWR _01912_ sky130_fd_sc_hd__mux2_1
XFILLER_0_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1013 _05468_ VGND VGND VPWR VPWR net1013 sky130_fd_sc_hd__buf_1
Xfanout1024 net1027 VGND VGND VPWR VPWR net1024 sky130_fd_sc_hd__clkbuf_2
XFILLER_126_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1035 _05458_ VGND VGND VPWR VPWR net1035 sky130_fd_sc_hd__buf_1
Xfanout1046 net1047 VGND VGND VPWR VPWR net1046 sky130_fd_sc_hd__clkbuf_2
Xfanout1057 _05446_ VGND VGND VPWR VPWR net1057 sky130_fd_sc_hd__clkbuf_1
X_10095_ net3081 net742 net638 VGND VGND VPWR VPWR _01844_ sky130_fd_sc_hd__mux2_1
Xfanout1068 _05440_ VGND VGND VPWR VPWR net1068 sky130_fd_sc_hd__clkbuf_2
Xfanout1079 _05436_ VGND VGND VPWR VPWR net1079 sky130_fd_sc_hd__clkbuf_2
X_13923_ clknet_leaf_220_clk _02552_ VGND VGND VPWR VPWR data_array.data1\[4\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_210_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_210_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_75_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13854_ clknet_leaf_24_clk _02483_ VGND VGND VPWR VPWR data_array.data1\[3\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12805_ clknet_leaf_130_clk _01499_ VGND VGND VPWR VPWR tag_array.tag1\[10\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_76_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13785_ clknet_leaf_254_clk _02414_ VGND VGND VPWR VPWR data_array.data1\[2\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_10997_ net1910 net1013 net341 VGND VGND VPWR VPWR _02741_ sky130_fd_sc_hd__mux2_1
XFILLER_31_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1036 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12736_ clknet_leaf_177_clk _01430_ VGND VGND VPWR VPWR tag_array.tag0\[5\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_700 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12667_ clknet_leaf_54_clk _01361_ VGND VGND VPWR VPWR data_array.data0\[15\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_61_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14406_ clknet_leaf_21_clk _03029_ VGND VGND VPWR VPWR data_array.data1\[10\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
X_11618_ clknet_leaf_127_clk _00426_ VGND VGND VPWR VPWR tag_array.tag1\[3\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_12598_ clknet_leaf_141_clk _01292_ VGND VGND VPWR VPWR tag_array.tag0\[0\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_14337_ clknet_leaf_238_clk _02966_ VGND VGND VPWR VPWR data_array.data1\[11\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
X_11549_ clknet_leaf_98_clk _00357_ VGND VGND VPWR VPWR tag_array.tag1\[6\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold507 data_array.data1\[8\]\[17\] VGND VGND VPWR VPWR net2158 sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 data_array.data0\[1\]\[5\] VGND VGND VPWR VPWR net2169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold529 data_array.data0\[4\]\[50\] VGND VGND VPWR VPWR net2180 sky130_fd_sc_hd__dlygate4sd3_1
X_14268_ clknet_leaf_210_clk _02897_ VGND VGND VPWR VPWR data_array.data1\[12\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_125_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13219_ clknet_leaf_12_clk _00115_ VGND VGND VPWR VPWR data_array.rdata1\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_131_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14199_ clknet_leaf_39_clk _02828_ VGND VGND VPWR VPWR data_array.data0\[2\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_111_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1207 data_array.data1\[13\]\[13\] VGND VGND VPWR VPWR net2858 sky130_fd_sc_hd__dlygate4sd3_1
X_08760_ net785 net3487 net450 VGND VGND VPWR VPWR _00519_ sky130_fd_sc_hd__mux2_1
XFILLER_140_997 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_05972_ data_array.rdata0\[47\] net1658 net1149 VGND VGND VPWR VPWR _03442_ sky130_fd_sc_hd__o21a_1
Xhold1218 data_array.data0\[9\]\[0\] VGND VGND VPWR VPWR net2869 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1229 tag_array.tag1\[2\]\[19\] VGND VGND VPWR VPWR net2880 sky130_fd_sc_hd__dlygate4sd3_1
X_07711_ data_array.data1\[1\]\[24\] net1578 net1482 data_array.data1\[2\]\[24\] VGND
+ VGND VPWR VPWR _04928_ sky130_fd_sc_hd__a22o_1
Xfanout1580 net1582 VGND VGND VPWR VPWR net1580 sky130_fd_sc_hd__clkbuf_4
Xfanout1591 _03508_ VGND VGND VPWR VPWR net1591 sky130_fd_sc_hd__buf_4
X_08691_ net2330 net760 net488 VGND VGND VPWR VPWR _00450_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_105_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_201_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_201_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07642_ data_array.data1\[4\]\[18\] net1345 net1251 data_array.data1\[7\]\[18\] _04864_
+ VGND VGND VPWR VPWR _04865_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_140_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07573_ data_array.data1\[9\]\[12\] net1586 net1490 data_array.data1\[10\]\[12\]
+ VGND VGND VPWR VPWR _04802_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_101_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09312_ net730 net2704 net548 VGND VGND VPWR VPWR _01066_ sky130_fd_sc_hd__mux2_1
X_06524_ tag_array.tag1\[4\]\[5\] net1420 net1326 tag_array.tag1\[7\]\[5\] _03848_
+ VGND VGND VPWR VPWR _03849_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_81_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09243_ net708 net2609 net646 VGND VGND VPWR VPWR _00997_ sky130_fd_sc_hd__mux2_1
XFILLER_166_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06455_ tag_array.tag0\[13\]\[24\] net1565 net1469 tag_array.tag0\[14\]\[24\] VGND
+ VGND VPWR VPWR _03786_ sky130_fd_sc_hd__a22o_1
XFILLER_21_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06386_ tag_array.tag0\[12\]\[18\] net1374 net1280 tag_array.tag0\[15\]\[18\] _03722_
+ VGND VGND VPWR VPWR _03723_ sky130_fd_sc_hd__a221o_1
X_09174_ net784 net3564 net627 VGND VGND VPWR VPWR _00928_ sky130_fd_sc_hd__mux2_1
XFILLER_147_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_268_clk clknet_5_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_268_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_175_872 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08125_ data_array.data1\[5\]\[62\] net1605 net1509 data_array.data1\[6\]\[62\] VGND
+ VGND VPWR VPWR _05304_ sky130_fd_sc_hd__a22o_1
XFILLER_147_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08056_ _05240_ _05241_ VGND VGND VPWR VPWR _00114_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_116_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07007_ data_array.data0\[1\]\[24\] net1577 net1481 data_array.data0\[2\]\[24\] VGND
+ VGND VPWR VPWR _04288_ sky130_fd_sc_hd__a22o_1
XFILLER_122_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_164_3515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput105 mem_rdata[15] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_1
Xinput116 mem_rdata[25] VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2420 tag_array.tag0\[0\]\[5\] VGND VGND VPWR VPWR net4071 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_181_3840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput127 mem_rdata[35] VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_1
Xhold2431 data_array.data0\[12\]\[16\] VGND VGND VPWR VPWR net4082 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput138 mem_rdata[45] VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_1
Xhold2442 tag_array.tag1\[10\]\[14\] VGND VGND VPWR VPWR net4093 sky130_fd_sc_hd__dlygate4sd3_1
X_08958_ net932 net4238 net432 VGND VGND VPWR VPWR _00714_ sky130_fd_sc_hd__mux2_1
Xinput149 mem_rdata[55] VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_1
Xhold2453 tag_array.tag0\[11\]\[23\] VGND VGND VPWR VPWR net4104 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2464 data_array.data0\[11\]\[47\] VGND VGND VPWR VPWR net4115 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1730 data_array.data1\[14\]\[25\] VGND VGND VPWR VPWR net3381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2475 data_array.data1\[6\]\[3\] VGND VGND VPWR VPWR net4126 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2486 data_array.data1\[10\]\[42\] VGND VGND VPWR VPWR net4137 sky130_fd_sc_hd__dlygate4sd3_1
X_07909_ data_array.data1\[1\]\[42\] net1585 net1489 data_array.data1\[2\]\[42\] VGND
+ VGND VPWR VPWR _05108_ sky130_fd_sc_hd__a22o_1
XFILLER_5_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1741 data_array.data0\[6\]\[24\] VGND VGND VPWR VPWR net3392 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1752 data_array.data1\[6\]\[53\] VGND VGND VPWR VPWR net3403 sky130_fd_sc_hd__dlygate4sd3_1
X_08889_ net948 net4260 net440 VGND VGND VPWR VPWR _00646_ sky130_fd_sc_hd__mux2_1
Xhold2497 data_array.data1\[5\]\[57\] VGND VGND VPWR VPWR net4148 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1763 data_array.data1\[5\]\[45\] VGND VGND VPWR VPWR net3414 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1774 tag_array.tag1\[6\]\[12\] VGND VGND VPWR VPWR net3425 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_5_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1785 tag_array.tag1\[9\]\[0\] VGND VGND VPWR VPWR net3436 sky130_fd_sc_hd__dlygate4sd3_1
X_10920_ net1062 net4620 net532 VGND VGND VPWR VPWR _02665_ sky130_fd_sc_hd__mux2_1
XFILLER_72_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1796 tag_array.tag0\[2\]\[13\] VGND VGND VPWR VPWR net3447 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_147_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10851_ net1082 net3711 net520 VGND VGND VPWR VPWR _02596_ sky130_fd_sc_hd__mux2_1
XFILLER_72_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_179_3791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13570_ clknet_leaf_28_clk _02199_ VGND VGND VPWR VPWR tag_array.dirty1\[4\] sky130_fd_sc_hd__dfxtp_1
X_10782_ net2002 net1100 net504 VGND VGND VPWR VPWR _02527_ sky130_fd_sc_hd__mux2_1
X_12521_ clknet_leaf_189_clk _01215_ VGND VGND VPWR VPWR tag_array.tag1\[11\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_23_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12452_ clknet_leaf_68_clk _01146_ VGND VGND VPWR VPWR data_array.data1\[9\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_36_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11403_ clknet_leaf_128_clk _00213_ VGND VGND VPWR VPWR tag_array.tag1\[7\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_259_clk clknet_5_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_259_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12383_ clknet_leaf_261_clk _01077_ VGND VGND VPWR VPWR data_array.data0\[14\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_14122_ clknet_leaf_11_clk _02751_ VGND VGND VPWR VPWR data_array.data0\[1\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11334_ net958 net4505 net802 VGND VGND VPWR VPWR _03077_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14053_ clknet_leaf_41_clk _02682_ VGND VGND VPWR VPWR data_array.data1\[6\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_11265_ net968 net3639 net673 VGND VGND VPWR VPWR _03008_ sky130_fd_sc_hd__mux2_1
XFILLER_180_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13004_ clknet_leaf_59_clk _01698_ VGND VGND VPWR VPWR data_array.data0\[3\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_122_942 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10216_ net940 net3351 net360 VGND VGND VPWR VPWR _01963_ sky130_fd_sc_hd__mux2_1
X_11196_ net991 net4207 net656 VGND VGND VPWR VPWR _02939_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10147_ net957 net3800 net366 VGND VGND VPWR VPWR _01895_ sky130_fd_sc_hd__mux2_1
XFILLER_79_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_85_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10078_ net713 net4182 net599 VGND VGND VPWR VPWR _01827_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_85_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13906_ clknet_leaf_115_clk _02535_ VGND VGND VPWR VPWR data_array.data1\[4\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13837_ clknet_leaf_198_clk _02466_ VGND VGND VPWR VPWR data_array.data1\[3\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_63_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13768_ clknet_leaf_227_clk _02397_ VGND VGND VPWR VPWR data_array.data1\[2\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_12719_ clknet_leaf_155_clk _01413_ VGND VGND VPWR VPWR tag_array.tag0\[7\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_13699_ clknet_leaf_41_clk _02328_ VGND VGND VPWR VPWR data_array.data1\[15\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_175_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06240_ net1174 _03585_ _03589_ net1221 VGND VGND VPWR VPWR _03591_ sky130_fd_sc_hd__a22o_1
XFILLER_176_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06171_ tag_array.valid0\[5\] net1597 net1501 tag_array.valid0\[6\] VGND VGND VPWR
+ VPWR _03528_ sky130_fd_sc_hd__a22o_1
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold304 data_array.data1\[5\]\[15\] VGND VGND VPWR VPWR net1955 sky130_fd_sc_hd__dlygate4sd3_1
Xhold315 data_array.data0\[5\]\[49\] VGND VGND VPWR VPWR net1966 sky130_fd_sc_hd__dlygate4sd3_1
Xhold326 data_array.data0\[4\]\[14\] VGND VGND VPWR VPWR net1977 sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 data_array.data0\[4\]\[7\] VGND VGND VPWR VPWR net1988 sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 data_array.data0\[1\]\[55\] VGND VGND VPWR VPWR net1999 sky130_fd_sc_hd__dlygate4sd3_1
X_09930_ net1108 net3554 net374 VGND VGND VPWR VPWR _01679_ sky130_fd_sc_hd__mux2_1
Xhold359 data_array.data1\[8\]\[12\] VGND VGND VPWR VPWR net2010 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout806 _05362_ VGND VGND VPWR VPWR net806 sky130_fd_sc_hd__buf_4
X_09861_ net1026 net2450 net380 VGND VGND VPWR VPWR _01611_ sky130_fd_sc_hd__mux2_1
Xfanout817 net818 VGND VGND VPWR VPWR net817 sky130_fd_sc_hd__clkbuf_4
XFILLER_124_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout828 net829 VGND VGND VPWR VPWR net828 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_74_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout839 net840 VGND VGND VPWR VPWR net839 sky130_fd_sc_hd__clkbuf_4
X_08812_ net2260 net998 net443 VGND VGND VPWR VPWR _00570_ sky130_fd_sc_hd__mux2_1
X_09792_ net1043 net3871 net386 VGND VGND VPWR VPWR _01543_ sky130_fd_sc_hd__mux2_1
Xhold1004 data_array.data0\[6\]\[49\] VGND VGND VPWR VPWR net2655 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1015 tag_array.tag0\[14\]\[7\] VGND VGND VPWR VPWR net2666 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_86_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1026 tag_array.tag0\[0\]\[19\] VGND VGND VPWR VPWR net2677 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1037 tag_array.tag0\[6\]\[6\] VGND VGND VPWR VPWR net2688 sky130_fd_sc_hd__dlygate4sd3_1
X_08743_ net750 net3173 net464 VGND VGND VPWR VPWR _00502_ sky130_fd_sc_hd__mux2_1
Xhold1048 data_array.data0\[8\]\[38\] VGND VGND VPWR VPWR net2699 sky130_fd_sc_hd__dlygate4sd3_1
X_05955_ data_array.rdata1\[41\] net829 net837 VGND VGND VPWR VPWR _03431_ sky130_fd_sc_hd__a21o_1
Xhold1059 data_array.data1\[11\]\[56\] VGND VGND VPWR VPWR net2710 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_54_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08674_ net728 net3634 net500 VGND VGND VPWR VPWR _00433_ sky130_fd_sc_hd__mux2_1
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05886_ data_array.rdata1\[18\] net829 net838 VGND VGND VPWR VPWR _03385_ sky130_fd_sc_hd__a21o_1
XFILLER_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07625_ net1621 _04843_ _04847_ net1195 VGND VGND VPWR VPWR _04850_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07556_ data_array.data1\[12\]\[10\] net1416 net1322 data_array.data1\[15\]\[10\]
+ _04786_ VGND VGND VPWR VPWR _04787_ sky130_fd_sc_hd__a221o_1
XFILLER_53_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06507_ tag_array.tag1\[8\]\[4\] net1362 net1268 tag_array.tag1\[11\]\[4\] _03832_
+ VGND VGND VPWR VPWR _03833_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_157_3374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07487_ data_array.data1\[5\]\[4\] net1583 net1487 data_array.data1\[6\]\[4\] VGND
+ VGND VPWR VPWR _04724_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_157_3385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09226_ net777 net2592 net645 VGND VGND VPWR VPWR _00980_ sky130_fd_sc_hd__mux2_1
X_06438_ net1174 _03765_ _03769_ net1221 VGND VGND VPWR VPWR _03771_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_118_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09157_ net914 net2817 net573 VGND VGND VPWR VPWR _00911_ sky130_fd_sc_hd__mux2_1
X_06369_ tag_array.tag0\[1\]\[16\] net1597 net1501 tag_array.tag0\[2\]\[16\] VGND
+ VGND VPWR VPWR _03708_ sky130_fd_sc_hd__a22o_1
XFILLER_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08108_ data_array.data1\[0\]\[60\] net1414 net1320 data_array.data1\[3\]\[60\] _05288_
+ VGND VGND VPWR VPWR _05289_ sky130_fd_sc_hd__a221o_1
XFILLER_181_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09088_ net932 net4112 net417 VGND VGND VPWR VPWR _00842_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_169_Right_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08039_ data_array.data1\[13\]\[54\] net1544 net1448 data_array.data1\[14\]\[54\]
+ VGND VGND VPWR VPWR _05226_ sky130_fd_sc_hd__a22o_1
XFILLER_107_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold860 tag_array.tag0\[0\]\[21\] VGND VGND VPWR VPWR net2511 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold871 data_array.data1\[12\]\[56\] VGND VGND VPWR VPWR net2522 sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 tag_array.tag0\[7\]\[23\] VGND VGND VPWR VPWR net2533 sky130_fd_sc_hd__dlygate4sd3_1
Xhold893 data_array.data1\[15\]\[14\] VGND VGND VPWR VPWR net2544 sky130_fd_sc_hd__dlygate4sd3_1
X_11050_ net2171 net1060 net335 VGND VGND VPWR VPWR _02793_ sky130_fd_sc_hd__mux2_1
XFILLER_27_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10001_ net1082 net2712 net563 VGND VGND VPWR VPWR _01750_ sky130_fd_sc_hd__mux2_1
XFILLER_153_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2250 data_array.data1\[6\]\[48\] VGND VGND VPWR VPWR net3901 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2261 data_array.data1\[13\]\[1\] VGND VGND VPWR VPWR net3912 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2272 tag_array.tag1\[10\]\[23\] VGND VGND VPWR VPWR net3923 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2283 data_array.data0\[14\]\[63\] VGND VGND VPWR VPWR net3934 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2294 tag_array.tag0\[7\]\[10\] VGND VGND VPWR VPWR net3945 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1560 tag_array.tag0\[6\]\[1\] VGND VGND VPWR VPWR net3211 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1571 data_array.data0\[3\]\[19\] VGND VGND VPWR VPWR net3222 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11952_ clknet_leaf_247_clk _00760_ VGND VGND VPWR VPWR data_array.data0\[4\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_28_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1582 data_array.data1\[12\]\[41\] VGND VGND VPWR VPWR net3233 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_28_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1593 tag_array.dirty1\[4\] VGND VGND VPWR VPWR net3244 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10903_ net875 net4504 net519 VGND VGND VPWR VPWR _02648_ sky130_fd_sc_hd__mux2_1
XFILLER_45_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11883_ clknet_leaf_228_clk _00691_ VGND VGND VPWR VPWR data_array.data0\[5\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_44_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13622_ clknet_leaf_38_clk _02251_ VGND VGND VPWR VPWR data_array.data0\[9\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
X_10834_ net2971 net892 net505 VGND VGND VPWR VPWR _02579_ sky130_fd_sc_hd__mux2_1
XFILLER_41_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13553_ clknet_leaf_246_clk _02182_ VGND VGND VPWR VPWR data_array.data1\[0\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_41_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10765_ net914 net4500 net497 VGND VGND VPWR VPWR _02510_ sky130_fd_sc_hd__mux2_1
XFILLER_157_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12504_ clknet_leaf_21_clk _01198_ VGND VGND VPWR VPWR data_array.data1\[9\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_158_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13484_ clknet_leaf_163_clk _02114_ VGND VGND VPWR VPWR tag_array.tag0\[15\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_121_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10696_ net2238 net934 net485 VGND VGND VPWR VPWR _02441_ sky130_fd_sc_hd__mux2_1
XFILLER_139_850 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12435_ clknet_leaf_3_clk _01129_ VGND VGND VPWR VPWR data_array.data0\[14\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12366_ clknet_leaf_76_clk _00042_ VGND VGND VPWR VPWR data_array.rdata0\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_136_Right_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14105_ clknet_leaf_249_clk _02734_ VGND VGND VPWR VPWR data_array.data0\[1\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_39_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11317_ net1024 net3188 net799 VGND VGND VPWR VPWR _03060_ sky130_fd_sc_hd__mux2_1
XFILLER_4_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12297_ clknet_leaf_195_clk _01055_ VGND VGND VPWR VPWR tag_array.tag1\[12\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_107_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_395 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14036_ clknet_leaf_86_clk _02665_ VGND VGND VPWR VPWR data_array.data1\[6\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_11248_ net1039 net4254 net675 VGND VGND VPWR VPWR _02991_ sky130_fd_sc_hd__mux2_1
XFILLER_80_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11179_ net1057 net3280 net652 VGND VGND VPWR VPWR _02922_ sky130_fd_sc_hd__mux2_1
XFILLER_67_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05740_ net5 fsm.tag_out1\[6\] VGND VGND VPWR VPWR _03257_ sky130_fd_sc_hd__and2b_1
XFILLER_169_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_704 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_05671_ net14 fsm.tag_out0\[14\] VGND VGND VPWR VPWR _03188_ sky130_fd_sc_hd__and2b_1
XFILLER_24_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07410_ data_array.data0\[1\]\[61\] net1548 net1452 data_array.data0\[2\]\[61\] VGND
+ VGND VPWR VPWR _04654_ sky130_fd_sc_hd__a22o_1
XFILLER_91_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08390_ net2418 net956 net691 VGND VGND VPWR VPWR _00259_ sky130_fd_sc_hd__mux2_1
XFILLER_149_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07341_ _04590_ _04591_ VGND VGND VPWR VPWR _00049_ sky130_fd_sc_hd__or2_1
XFILLER_177_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07272_ data_array.data0\[0\]\[48\] net1381 net1287 data_array.data0\[3\]\[48\] _04528_
+ VGND VGND VPWR VPWR _04529_ sky130_fd_sc_hd__a221o_1
XFILLER_177_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09011_ net2016 net982 net418 VGND VGND VPWR VPWR _00766_ sky130_fd_sc_hd__mux2_1
XFILLER_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06223_ tag_array.tag0\[0\]\[3\] net1371 net1277 tag_array.tag0\[3\]\[3\] _03574_
+ VGND VGND VPWR VPWR _03575_ sky130_fd_sc_hd__a221o_1
XFILLER_163_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06154_ net26 net27 VGND VGND VPWR VPWR _03511_ sky130_fd_sc_hd__nand2b_2
XFILLER_129_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold101 data_array.data0\[1\]\[25\] VGND VGND VPWR VPWR net1752 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold112 data_array.data0\[2\]\[62\] VGND VGND VPWR VPWR net1763 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 data_array.data1\[0\]\[26\] VGND VGND VPWR VPWR net1774 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold134 data_array.data1\[0\]\[17\] VGND VGND VPWR VPWR net1785 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_103_Right_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06085_ data_array.rdata0\[0\] net1137 net1118 data_array.rdata1\[0\] VGND VGND VPWR
+ VPWR net263 sky130_fd_sc_hd__a22o_1
Xhold145 data_array.data1\[8\]\[11\] VGND VGND VPWR VPWR net1796 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold156 tag_array.tag1\[0\]\[0\] VGND VGND VPWR VPWR net1807 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 data_array.data1\[4\]\[19\] VGND VGND VPWR VPWR net1818 sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 data_array.data1\[0\]\[2\] VGND VGND VPWR VPWR net1829 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_99_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09913_ net754 net2941 net603 VGND VGND VPWR VPWR _01663_ sky130_fd_sc_hd__mux2_1
Xfanout603 net604 VGND VGND VPWR VPWR net603 sky130_fd_sc_hd__buf_4
Xhold189 tag_array.tag1\[0\]\[19\] VGND VGND VPWR VPWR net1840 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout614 _05573_ VGND VGND VPWR VPWR net614 sky130_fd_sc_hd__buf_4
Xfanout625 _05565_ VGND VGND VPWR VPWR net625 sky130_fd_sc_hd__buf_4
Xfanout636 _05557_ VGND VGND VPWR VPWR net636 sky130_fd_sc_hd__clkbuf_4
X_09844_ net1093 net3347 net383 VGND VGND VPWR VPWR _01594_ sky130_fd_sc_hd__mux2_1
Xfanout647 _05555_ VGND VGND VPWR VPWR net647 sky130_fd_sc_hd__buf_4
Xfanout658 net659 VGND VGND VPWR VPWR net658 sky130_fd_sc_hd__buf_4
XFILLER_58_336 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout669 net670 VGND VGND VPWR VPWR net669 sky130_fd_sc_hd__buf_2
XFILLER_37_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09775_ net1109 net3105 net389 VGND VGND VPWR VPWR _01526_ sky130_fd_sc_hd__mux2_1
X_06987_ net1618 _04263_ _04267_ net1192 VGND VGND VPWR VPWR _04270_ sky130_fd_sc_hd__a22o_1
XFILLER_39_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08726_ net1732 net718 net470 VGND VGND VPWR VPWR _00485_ sky130_fd_sc_hd__mux2_1
XFILLER_113_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05938_ net127 net1150 _03418_ _03419_ VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__a22o_1
XFILLER_2_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_3414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08657_ net2648 net694 net506 VGND VGND VPWR VPWR _00416_ sky130_fd_sc_hd__mux2_1
X_05869_ net102 net1157 _03372_ _03373_ VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__a22o_1
XFILLER_163_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_3425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07608_ data_array.data1\[5\]\[15\] net1584 net1488 data_array.data1\[6\]\[15\] VGND
+ VGND VPWR VPWR _04834_ sky130_fd_sc_hd__a22o_1
X_08588_ net773 net3944 net535 VGND VGND VPWR VPWR _00347_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_176_3750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07539_ _04770_ _04771_ VGND VGND VPWR VPWR _00126_ sky130_fd_sc_hd__or2_1
XFILLER_23_984 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10550_ net1004 net3503 net454 VGND VGND VPWR VPWR _02295_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_172_3669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09209_ net744 net2848 net630 VGND VGND VPWR VPWR _00963_ sky130_fd_sc_hd__mux2_1
XFILLER_33_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10481_ net1022 net3681 net345 VGND VGND VPWR VPWR _02226_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_133_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12220_ clknet_leaf_151_clk _00173_ VGND VGND VPWR VPWR fsm.tag_out1\[2\] sky130_fd_sc_hd__dfxtp_1
X_12151_ clknet_leaf_145_clk _00959_ VGND VGND VPWR VPWR tag_array.tag0\[13\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_162_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11102_ net1111 net3770 net546 VGND VGND VPWR VPWR _02845_ sky130_fd_sc_hd__mux2_1
XFILLER_123_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12082_ clknet_leaf_30_clk _00890_ VGND VGND VPWR VPWR data_array.data1\[14\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_111_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold690 data_array.data0\[10\]\[52\] VGND VGND VPWR VPWR net2341 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11033_ net2436 net868 net343 VGND VGND VPWR VPWR _02777_ sky130_fd_sc_hd__mux2_1
XFILLER_104_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2080 data_array.data1\[14\]\[18\] VGND VGND VPWR VPWR net3731 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2091 data_array.data0\[13\]\[57\] VGND VGND VPWR VPWR net3742 sky130_fd_sc_hd__dlygate4sd3_1
X_12984_ clknet_leaf_186_clk _01678_ VGND VGND VPWR VPWR tag_array.tag0\[4\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1390 data_array.data0\[3\]\[13\] VGND VGND VPWR VPWR net3041 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11935_ clknet_leaf_62_clk _00743_ VGND VGND VPWR VPWR data_array.data0\[4\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11866_ clknet_leaf_72_clk _00674_ VGND VGND VPWR VPWR data_array.data0\[5\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_13605_ clknet_leaf_70_clk _02234_ VGND VGND VPWR VPWR data_array.data0\[9\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_10817_ net1986 net960 net505 VGND VGND VPWR VPWR _02562_ sky130_fd_sc_hd__mux2_1
X_11797_ clknet_leaf_224_clk _00605_ VGND VGND VPWR VPWR data_array.data0\[8\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13536_ clknet_leaf_73_clk _02165_ VGND VGND VPWR VPWR data_array.data1\[0\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
X_10748_ net980 net3710 net490 VGND VGND VPWR VPWR _02493_ sky130_fd_sc_hd__mux2_1
XFILLER_146_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13467_ clknet_leaf_108_clk _02097_ VGND VGND VPWR VPWR tag_array.tag0\[1\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_146_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10679_ net2025 net1000 net478 VGND VGND VPWR VPWR _02424_ sky130_fd_sc_hd__mux2_1
XFILLER_173_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12418_ clknet_leaf_85_clk _01112_ VGND VGND VPWR VPWR data_array.data0\[14\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_127_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13398_ clknet_leaf_19_clk _02028_ VGND VGND VPWR VPWR data_array.data1\[8\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput206 net206 VGND VGND VPWR VPWR cpu_rdata[47] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_93_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput217 net217 VGND VGND VPWR VPWR cpu_rdata[57] sky130_fd_sc_hd__clkbuf_4
XFILLER_126_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput228 net228 VGND VGND VPWR VPWR cpu_rdata[9] sky130_fd_sc_hd__buf_6
XFILLER_5_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12349_ clknet_leaf_49_clk _00024_ VGND VGND VPWR VPWR data_array.rdata0\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_154_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput239 net239 VGND VGND VPWR VPWR mem_addr[18] sky130_fd_sc_hd__buf_2
XFILLER_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06910_ net1632 _04193_ _04197_ net1206 VGND VGND VPWR VPWR _04200_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_71_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14019_ clknet_leaf_54_clk _02648_ VGND VGND VPWR VPWR data_array.data1\[5\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07890_ net1185 _05085_ _05089_ net1231 VGND VGND VPWR VPWR _05091_ sky130_fd_sc_hd__a22o_1
XFILLER_68_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06841_ data_array.data0\[12\]\[9\] net1389 net1295 data_array.data0\[15\]\[9\] _04136_
+ VGND VGND VPWR VPWR _04137_ sky130_fd_sc_hd__a221o_1
XFILLER_95_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09560_ net1109 net4061 net397 VGND VGND VPWR VPWR _01312_ sky130_fd_sc_hd__mux2_1
XFILLER_110_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06772_ data_array.data0\[5\]\[3\] net1567 net1471 data_array.data0\[6\]\[3\] VGND
+ VGND VPWR VPWR _04074_ sky130_fd_sc_hd__a22o_1
X_08511_ _03509_ _03527_ net821 VGND VGND VPWR VPWR _05578_ sky130_fd_sc_hd__or3_1
X_05723_ net3 fsm.tag_out1\[4\] VGND VGND VPWR VPWR _03240_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_19_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09491_ net762 net4408 net626 VGND VGND VPWR VPWR _01244_ sky130_fd_sc_hd__mux2_1
XFILLER_64_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08442_ net150 net85 net1639 VGND VGND VPWR VPWR _05531_ sky130_fd_sc_hd__mux2_1
X_05654_ _03167_ _03168_ _03169_ _03170_ VGND VGND VPWR VPWR _03171_ sky130_fd_sc_hd__or4_1
XFILLER_23_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08373_ net125 net60 net1641 VGND VGND VPWR VPWR _05485_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_154_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07324_ data_array.data0\[13\]\[53\] net1522 net1426 data_array.data0\[14\]\[53\]
+ VGND VGND VPWR VPWR _04576_ sky130_fd_sc_hd__a22o_1
XFILLER_104_1004 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07255_ data_array.data0\[8\]\[47\] net1387 net1293 data_array.data0\[11\]\[47\]
+ _04512_ VGND VGND VPWR VPWR _04513_ sky130_fd_sc_hd__a221o_1
XFILLER_176_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06206_ net1633 _03553_ _03557_ net1207 VGND VGND VPWR VPWR _03560_ sky130_fd_sc_hd__a22o_1
XFILLER_136_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07186_ net1183 _04445_ _04449_ net1231 VGND VGND VPWR VPWR _04451_ sky130_fd_sc_hd__a22o_1
XFILLER_173_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06137_ data_array.rdata0\[52\] net1136 net1117 data_array.rdata1\[52\] VGND VGND
+ VPWR VPWR net310 sky130_fd_sc_hd__a22o_1
XFILLER_133_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06068_ fsm.tag_out0\[16\] net1121 _03497_ VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__a21o_1
Xfanout400 net401 VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__clkbuf_8
Xfanout411 net417 VGND VGND VPWR VPWR net411 sky130_fd_sc_hd__clkbuf_4
Xfanout1409 net1422 VGND VGND VPWR VPWR net1409 sky130_fd_sc_hd__clkbuf_4
XFILLER_87_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout422 net423 VGND VGND VPWR VPWR net422 sky130_fd_sc_hd__buf_4
Xfanout433 _05609_ VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__buf_6
XFILLER_58_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout444 net445 VGND VGND VPWR VPWR net444 sky130_fd_sc_hd__buf_4
XFILLER_58_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout455 net459 VGND VGND VPWR VPWR net455 sky130_fd_sc_hd__clkbuf_8
XFILLER_113_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout466 net468 VGND VGND VPWR VPWR net466 sky130_fd_sc_hd__clkbuf_8
XFILLER_87_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09827_ net903 net4142 net388 VGND VGND VPWR VPWR _01578_ sky130_fd_sc_hd__mux2_1
Xfanout477 _05603_ VGND VGND VPWR VPWR net477 sky130_fd_sc_hd__clkbuf_4
XFILLER_74_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout488 net489 VGND VGND VPWR VPWR net488 sky130_fd_sc_hd__buf_4
XFILLER_74_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout499 _05601_ VGND VGND VPWR VPWR net499 sky130_fd_sc_hd__buf_4
X_09758_ net3693 net756 net671 VGND VGND VPWR VPWR _01510_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_126_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08709_ net1784 net787 net471 VGND VGND VPWR VPWR _00468_ sky130_fd_sc_hd__mux2_1
X_09689_ net732 net3974 net606 VGND VGND VPWR VPWR _01441_ sky130_fd_sc_hd__mux2_1
XFILLER_27_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11720_ clknet_leaf_165_clk _00528_ VGND VGND VPWR VPWR tag_array.tag0\[9\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_174_3709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11651_ clknet_leaf_128_clk _00459_ VGND VGND VPWR VPWR tag_array.tag1\[2\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10602_ net2262 net1054 net471 VGND VGND VPWR VPWR _02347_ sky130_fd_sc_hd__mux2_1
X_14370_ clknet_leaf_122_clk _02993_ VGND VGND VPWR VPWR data_array.data1\[10\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_11582_ clknet_leaf_129_clk _00390_ VGND VGND VPWR VPWR tag_array.tag1\[5\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_167_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13321_ clknet_leaf_70_clk _01951_ VGND VGND VPWR VPWR data_array.data0\[10\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_10533_ net1074 net4593 net461 VGND VGND VPWR VPWR _02278_ sky130_fd_sc_hd__mux2_1
XFILLER_167_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire845 _03236_ VGND VGND VPWR VPWR net845 sky130_fd_sc_hd__buf_2
XFILLER_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13252_ clknet_leaf_4_clk _01882_ VGND VGND VPWR VPWR data_array.data0\[11\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_10464_ net1089 net2421 net346 VGND VGND VPWR VPWR _02209_ sky130_fd_sc_hd__mux2_1
XFILLER_143_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12203_ clknet_leaf_145_clk _00132_ VGND VGND VPWR VPWR fsm.tag_out0\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_109_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13183_ clknet_leaf_122_clk _00076_ VGND VGND VPWR VPWR data_array.rdata1\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_136_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10395_ net2190 net1074 net668 VGND VGND VPWR VPWR _02141_ sky130_fd_sc_hd__mux2_1
XFILLER_151_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12134_ clknet_leaf_145_clk _00942_ VGND VGND VPWR VPWR tag_array.tag0\[12\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12065_ clknet_leaf_35_clk _00873_ VGND VGND VPWR VPWR data_array.data1\[14\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_111_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11016_ net2429 net936 net342 VGND VGND VPWR VPWR _02760_ sky130_fd_sc_hd__mux2_1
XFILLER_65_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_24__f_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_5_24__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_18_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12967_ clknet_leaf_143_clk _01661_ VGND VGND VPWR VPWR tag_array.tag0\[4\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_16_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11918_ clknet_leaf_12_clk _00726_ VGND VGND VPWR VPWR data_array.data0\[5\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_178_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12898_ clknet_leaf_247_clk _01592_ VGND VGND VPWR VPWR data_array.data0\[13\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_61_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11849_ clknet_leaf_1_clk _00657_ VGND VGND VPWR VPWR data_array.data0\[7\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13519_ clknet_leaf_214_clk _02148_ VGND VGND VPWR VPWR data_array.data1\[0\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_146_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14499_ clknet_leaf_181_clk _00128_ VGND VGND VPWR VPWR fsm.lru_out sky130_fd_sc_hd__dfxtp_1
Xclkload10 clknet_5_22__leaf_clk VGND VGND VPWR VPWR clkload10/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload21 clknet_leaf_6_clk VGND VGND VPWR VPWR clkload21/Y sky130_fd_sc_hd__inv_8
X_07040_ data_array.data0\[5\]\[27\] net1555 net1459 data_array.data0\[6\]\[27\] VGND
+ VGND VPWR VPWR _04318_ sky130_fd_sc_hd__a22o_1
XFILLER_146_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload32 clknet_leaf_12_clk VGND VGND VPWR VPWR clkload32/X sky130_fd_sc_hd__clkbuf_4
Xclkload43 clknet_leaf_23_clk VGND VGND VPWR VPWR clkload43/Y sky130_fd_sc_hd__inv_6
Xclkload54 clknet_leaf_252_clk VGND VGND VPWR VPWR clkload54/Y sky130_fd_sc_hd__inv_6
Xclkload65 clknet_leaf_243_clk VGND VGND VPWR VPWR clkload65/Y sky130_fd_sc_hd__inv_6
Xclkload76 clknet_leaf_48_clk VGND VGND VPWR VPWR clkload76/Y sky130_fd_sc_hd__clkinv_2
Xclkload87 clknet_leaf_55_clk VGND VGND VPWR VPWR clkload87/X sky130_fd_sc_hd__clkbuf_8
XFILLER_114_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload98 clknet_leaf_68_clk VGND VGND VPWR VPWR clkload98/Y sky130_fd_sc_hd__bufinv_16
XFILLER_86_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08991_ net2134 net1060 net424 VGND VGND VPWR VPWR _00746_ sky130_fd_sc_hd__mux2_1
XFILLER_141_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_1046 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2805 tag_array.tag1\[7\]\[12\] VGND VGND VPWR VPWR net4456 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2816 data_array.data0\[13\]\[23\] VGND VGND VPWR VPWR net4467 sky130_fd_sc_hd__dlygate4sd3_1
X_07942_ data_array.data1\[5\]\[45\] net1540 net1444 data_array.data1\[6\]\[45\] VGND
+ VGND VPWR VPWR _05138_ sky130_fd_sc_hd__a22o_1
Xhold2827 data_array.data1\[3\]\[17\] VGND VGND VPWR VPWR net4478 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_141_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2838 data_array.data1\[3\]\[1\] VGND VGND VPWR VPWR net4489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2849 data_array.data1\[3\]\[49\] VGND VGND VPWR VPWR net4500 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_147_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07873_ data_array.data1\[0\]\[39\] net1347 net1253 data_array.data1\[3\]\[39\] _05074_
+ VGND VGND VPWR VPWR _05075_ sky130_fd_sc_hd__a221o_1
XFILLER_96_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09612_ net903 net3550 net396 VGND VGND VPWR VPWR _01364_ sky130_fd_sc_hd__mux2_1
XFILLER_110_572 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_108_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06824_ _04120_ _04121_ VGND VGND VPWR VPWR _00061_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_108_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09543_ net754 net3134 net619 VGND VGND VPWR VPWR _01296_ sky130_fd_sc_hd__mux2_1
X_06755_ data_array.data0\[4\]\[1\] net1331 net1237 data_array.data0\[7\]\[1\] _04058_
+ VGND VGND VPWR VPWR _04059_ sky130_fd_sc_hd__a221o_1
XFILLER_36_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_05706_ _03163_ _03183_ _03201_ VGND VGND VPWR VPWR _03223_ sky130_fd_sc_hd__or3_1
X_09474_ net731 net3547 net655 VGND VGND VPWR VPWR _01227_ sky130_fd_sc_hd__mux2_1
X_06686_ tag_array.tag1\[13\]\[20\] net1558 net1462 tag_array.tag1\[14\]\[20\] VGND
+ VGND VPWR VPWR _03996_ sky130_fd_sc_hd__a22o_1
XFILLER_180_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08425_ net1123 _05519_ VGND VGND VPWR VPWR _05520_ sky130_fd_sc_hd__and2_1
X_05637_ fsm.state\[2\] net33 VGND VGND VPWR VPWR _03154_ sky130_fd_sc_hd__and2_4
XTAP_TAPCELL_ROW_121_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08356_ net1125 _05473_ VGND VGND VPWR VPWR _05474_ sky130_fd_sc_hd__and2_1
XFILLER_177_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload4 clknet_5_8__leaf_clk VGND VGND VPWR VPWR clkload4/X sky130_fd_sc_hd__clkbuf_8
X_07307_ net1167 _04555_ _04559_ net1213 VGND VGND VPWR VPWR _04561_ sky130_fd_sc_hd__a22o_1
XFILLER_50_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08287_ net1127 _05427_ VGND VGND VPWR VPWR _05428_ sky130_fd_sc_hd__and2_1
XFILLER_166_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07238_ data_array.data0\[5\]\[45\] net1535 net1439 data_array.data0\[6\]\[45\] VGND
+ VGND VPWR VPWR _04498_ sky130_fd_sc_hd__a22o_1
XFILLER_4_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07169_ data_array.data0\[0\]\[39\] net1348 net1254 data_array.data0\[3\]\[39\] _04434_
+ VGND VGND VPWR VPWR _04435_ sky130_fd_sc_hd__a221o_1
XFILLER_59_24 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10180_ net1084 net4271 net354 VGND VGND VPWR VPWR _01927_ sky130_fd_sc_hd__mux2_1
XFILLER_121_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_167_3568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_3579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1206 net1212 VGND VGND VPWR VPWR net1206 sky130_fd_sc_hd__buf_4
Xfanout1217 net1223 VGND VGND VPWR VPWR net1217 sky130_fd_sc_hd__buf_4
Xfanout1228 net1234 VGND VGND VPWR VPWR net1228 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_184_3893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1239 net1240 VGND VGND VPWR VPWR net1239 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_128_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13870_ clknet_leaf_74_clk _02499_ VGND VGND VPWR VPWR data_array.data1\[3\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_101_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12821_ clknet_leaf_168_clk _01515_ VGND VGND VPWR VPWR tag_array.tag1\[0\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12752_ clknet_leaf_169_clk _01446_ VGND VGND VPWR VPWR tag_array.tag0\[5\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_11703_ clknet_leaf_103_clk _00511_ VGND VGND VPWR VPWR tag_array.tag1\[15\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_12683_ clknet_leaf_163_clk _01377_ VGND VGND VPWR VPWR tag_array.tag0\[8\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_14422_ clknet_leaf_269_clk _03045_ VGND VGND VPWR VPWR data_array.data1\[7\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_91_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11634_ clknet_leaf_97_clk _00442_ VGND VGND VPWR VPWR tag_array.tag1\[2\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_156_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14353_ clknet_leaf_19_clk _02976_ VGND VGND VPWR VPWR data_array.data1\[10\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_156_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11565_ clknet_leaf_193_clk _00373_ VGND VGND VPWR VPWR tag_array.tag1\[5\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13304_ clknet_leaf_206_clk _01934_ VGND VGND VPWR VPWR data_array.data0\[10\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_42_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_907 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10516_ net880 net4150 net347 VGND VGND VPWR VPWR _02261_ sky130_fd_sc_hd__mux2_1
X_14284_ clknet_leaf_68_clk _02913_ VGND VGND VPWR VPWR data_array.data1\[11\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_21_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11496_ clknet_leaf_183_clk _00182_ VGND VGND VPWR VPWR fsm.valid1 sky130_fd_sc_hd__dfxtp_1
XFILLER_6_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13235_ clknet_leaf_16_clk _01865_ VGND VGND VPWR VPWR data_array.data0\[11\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_90_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10447_ net1851 net865 net665 VGND VGND VPWR VPWR _02193_ sky130_fd_sc_hd__mux2_1
XFILLER_3_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13166_ clknet_leaf_48_clk _00097_ VGND VGND VPWR VPWR data_array.rdata1\[3\] sky130_fd_sc_hd__dfxtp_1
X_10378_ net352 net2862 net580 VGND VGND VPWR VPWR _02124_ sky130_fd_sc_hd__mux2_1
X_12117_ clknet_leaf_192_clk _00925_ VGND VGND VPWR VPWR data_array.data1\[14\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13097_ clknet_leaf_75_clk _01791_ VGND VGND VPWR VPWR data_array.data1\[13\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_111_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12048_ clknet_leaf_208_clk _00856_ VGND VGND VPWR VPWR data_array.data0\[6\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_88_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_968 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13999_ clknet_leaf_236_clk _02628_ VGND VGND VPWR VPWR data_array.data1\[5\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
X_06540_ tag_array.tag1\[8\]\[7\] net1421 net1327 tag_array.tag1\[11\]\[7\] _03862_
+ VGND VGND VPWR VPWR _03863_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_66_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06471_ net1225 _03795_ _03799_ net1177 VGND VGND VPWR VPWR _03801_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_83_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08210_ fsm.tag_out1\[5\] net817 net809 net1653 _05374_ VGND VGND VPWR VPWR _05375_
+ sky130_fd_sc_hd__a221o_1
XFILLER_53_1031 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09190_ net720 net3546 net627 VGND VGND VPWR VPWR _00944_ sky130_fd_sc_hd__mux2_1
XFILLER_60_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08141_ data_array.data1\[0\]\[63\] net1361 net1267 data_array.data1\[3\]\[63\] _05318_
+ VGND VGND VPWR VPWR _05319_ sky130_fd_sc_hd__a221o_1
XFILLER_14_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08072_ data_array.data1\[9\]\[57\] net1538 net1442 data_array.data1\[10\]\[57\]
+ VGND VGND VPWR VPWR _05256_ sky130_fd_sc_hd__a22o_1
Xclkload110 clknet_leaf_93_clk VGND VGND VPWR VPWR clkload110/X sky130_fd_sc_hd__clkbuf_8
Xclkload121 clknet_leaf_88_clk VGND VGND VPWR VPWR clkload121/Y sky130_fd_sc_hd__clkinv_2
XFILLER_174_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload132 clknet_leaf_213_clk VGND VGND VPWR VPWR clkload132/Y sky130_fd_sc_hd__clkinv_4
Xclkload143 clknet_leaf_208_clk VGND VGND VPWR VPWR clkload143/Y sky130_fd_sc_hd__inv_6
XFILLER_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07023_ data_array.data0\[9\]\[26\] net1527 net1431 data_array.data0\[10\]\[26\]
+ VGND VGND VPWR VPWR _04302_ sky130_fd_sc_hd__a22o_1
Xclkload154 clknet_leaf_231_clk VGND VGND VPWR VPWR clkload154/Y sky130_fd_sc_hd__inv_6
XFILLER_161_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload165 clknet_leaf_203_clk VGND VGND VPWR VPWR clkload165/Y sky130_fd_sc_hd__clkinv_2
Xclkload176 clknet_leaf_176_clk VGND VGND VPWR VPWR clkload176/Y sky130_fd_sc_hd__clkinv_4
Xclkload187 clknet_leaf_188_clk VGND VGND VPWR VPWR clkload187/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_149_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload198 clknet_leaf_107_clk VGND VGND VPWR VPWR clkload198/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_149_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08974_ net869 net3463 net432 VGND VGND VPWR VPWR _00730_ sky130_fd_sc_hd__mux2_1
Xhold2602 data_array.data1\[15\]\[50\] VGND VGND VPWR VPWR net4253 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2613 data_array.data0\[13\]\[32\] VGND VGND VPWR VPWR net4264 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2624 data_array.data1\[3\]\[48\] VGND VGND VPWR VPWR net4275 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2635 data_array.data0\[14\]\[55\] VGND VGND VPWR VPWR net4286 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_89_Right_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07925_ data_array.data1\[9\]\[44\] net1590 net1494 data_array.data1\[10\]\[44\]
+ VGND VGND VPWR VPWR _05122_ sky130_fd_sc_hd__a22o_1
Xhold1901 tag_array.tag0\[9\]\[0\] VGND VGND VPWR VPWR net3552 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2646 data_array.data0\[6\]\[11\] VGND VGND VPWR VPWR net4297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2657 data_array.data1\[15\]\[46\] VGND VGND VPWR VPWR net4308 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_68_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold49 tag_array.valid1\[9\] VGND VGND VPWR VPWR net1700 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1912 data_array.data1\[3\]\[55\] VGND VGND VPWR VPWR net3563 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2668 data_array.data0\[9\]\[21\] VGND VGND VPWR VPWR net4319 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_68_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1923 tag_array.tag0\[6\]\[9\] VGND VGND VPWR VPWR net3574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2679 data_array.data0\[10\]\[34\] VGND VGND VPWR VPWR net4330 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1934 tag_array.tag0\[5\]\[12\] VGND VGND VPWR VPWR net3585 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_162_3476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1945 tag_array.tag0\[13\]\[1\] VGND VGND VPWR VPWR net3596 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1956 data_array.data0\[7\]\[5\] VGND VGND VPWR VPWR net3607 sky130_fd_sc_hd__dlygate4sd3_1
X_07856_ net1621 _05053_ _05057_ net1195 VGND VGND VPWR VPWR _05060_ sky130_fd_sc_hd__a22o_1
XFILLER_110_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1967 data_array.data0\[7\]\[61\] VGND VGND VPWR VPWR net3618 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1978 tag_array.tag0\[1\]\[16\] VGND VGND VPWR VPWR net3629 sky130_fd_sc_hd__dlygate4sd3_1
X_06807_ data_array.data0\[13\]\[6\] net1519 net1423 data_array.data0\[14\]\[6\] VGND
+ VGND VPWR VPWR _04106_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_123_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1989 data_array.data0\[7\]\[47\] VGND VGND VPWR VPWR net3640 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_16_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07787_ data_array.data1\[8\]\[31\] net1384 net1290 data_array.data1\[11\]\[31\]
+ _04996_ VGND VGND VPWR VPWR _04997_ sky130_fd_sc_hd__a221o_1
XFILLER_25_810 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09526_ net723 net3521 net622 VGND VGND VPWR VPWR _01279_ sky130_fd_sc_hd__mux2_1
X_06738_ data_array.data0\[12\]\[0\] net1365 net1271 data_array.data0\[15\]\[0\] _04042_
+ VGND VGND VPWR VPWR _04043_ sky130_fd_sc_hd__a221o_1
XFILLER_169_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09457_ net819 net3962 _05588_ VGND VGND VPWR VPWR _01210_ sky130_fd_sc_hd__mux2_1
X_06669_ net1221 _03975_ _03979_ net1172 VGND VGND VPWR VPWR _03981_ sky130_fd_sc_hd__a22o_1
XFILLER_80_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08408_ net2623 net932 _05417_ VGND VGND VPWR VPWR _00265_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_98_Right_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09388_ net819 net3404 _05572_ VGND VGND VPWR VPWR _01141_ sky130_fd_sc_hd__mux2_1
XFILLER_138_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08339_ net1825 net1027 net688 VGND VGND VPWR VPWR _00242_ sky130_fd_sc_hd__mux2_1
XFILLER_177_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11350_ net892 net4403 net798 VGND VGND VPWR VPWR _03093_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_169_3608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10301_ net3466 net958 net640 VGND VGND VPWR VPWR _02048_ sky130_fd_sc_hd__mux2_1
XFILLER_165_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11281_ net907 net3560 net673 VGND VGND VPWR VPWR _03024_ sky130_fd_sc_hd__mux2_1
XFILLER_137_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13020_ clknet_leaf_244_clk _01714_ VGND VGND VPWR VPWR data_array.data0\[3\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
X_10232_ net876 net3924 net356 VGND VGND VPWR VPWR _01979_ sky130_fd_sc_hd__mux2_1
XFILLER_180_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10163_ net894 net3712 net364 VGND VGND VPWR VPWR _01911_ sky130_fd_sc_hd__mux2_1
Xfanout1003 _05474_ VGND VGND VPWR VPWR net1003 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1014 net1015 VGND VGND VPWR VPWR net1014 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1025 net1027 VGND VGND VPWR VPWR net1025 sky130_fd_sc_hd__clkbuf_2
Xfanout1036 _05456_ VGND VGND VPWR VPWR net1036 sky130_fd_sc_hd__clkbuf_2
Xfanout1047 _05452_ VGND VGND VPWR VPWR net1047 sky130_fd_sc_hd__dlymetal6s2s_1
X_10094_ net1863 net747 net639 VGND VGND VPWR VPWR _01843_ sky130_fd_sc_hd__mux2_1
Xfanout1058 _05446_ VGND VGND VPWR VPWR net1058 sky130_fd_sc_hd__clkbuf_2
Xfanout1069 _05440_ VGND VGND VPWR VPWR net1069 sky130_fd_sc_hd__buf_1
X_13922_ clknet_leaf_254_clk _02551_ VGND VGND VPWR VPWR data_array.data1\[4\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_48_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_467 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13853_ clknet_leaf_228_clk _02482_ VGND VGND VPWR VPWR data_array.data1\[3\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_142_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12804_ clknet_leaf_197_clk _01498_ VGND VGND VPWR VPWR tag_array.tag1\[10\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_13784_ clknet_leaf_214_clk _02413_ VGND VGND VPWR VPWR data_array.data1\[2\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_10996_ net2303 net1018 net338 VGND VGND VPWR VPWR _02740_ sky130_fd_sc_hd__mux2_1
XFILLER_15_353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12735_ clknet_leaf_177_clk _01429_ VGND VGND VPWR VPWR tag_array.tag0\[5\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1048 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ clknet_leaf_57_clk _01360_ VGND VGND VPWR VPWR data_array.data0\[15\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_61_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_712 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14405_ clknet_leaf_17_clk _03028_ VGND VGND VPWR VPWR data_array.data1\[10\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
X_11617_ clknet_leaf_138_clk _00425_ VGND VGND VPWR VPWR tag_array.tag1\[3\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_12597_ clknet_leaf_177_clk _01291_ VGND VGND VPWR VPWR tag_array.tag0\[0\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_14336_ clknet_leaf_21_clk _02965_ VGND VGND VPWR VPWR data_array.data1\[11\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
X_11548_ clknet_leaf_232_clk _00356_ VGND VGND VPWR VPWR tag_array.tag1\[6\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold508 data_array.data1\[1\]\[61\] VGND VGND VPWR VPWR net2159 sky130_fd_sc_hd__dlygate4sd3_1
X_14267_ clknet_leaf_4_clk _02896_ VGND VGND VPWR VPWR data_array.data1\[12\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold519 data_array.data1\[13\]\[17\] VGND VGND VPWR VPWR net2170 sky130_fd_sc_hd__dlygate4sd3_1
X_11479_ clknet_leaf_156_clk _00288_ VGND VGND VPWR VPWR tag_array.valid0\[14\] sky130_fd_sc_hd__dfxtp_1
X_13218_ clknet_leaf_14_clk _00114_ VGND VGND VPWR VPWR data_array.rdata1\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_100_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14198_ clknet_leaf_6_clk _02827_ VGND VGND VPWR VPWR data_array.data0\[2\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_124_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13149_ clknet_leaf_32_clk _01843_ VGND VGND VPWR VPWR tag_array.tag1\[8\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1208 data_array.data0\[1\]\[20\] VGND VGND VPWR VPWR net2859 sky130_fd_sc_hd__dlygate4sd3_1
X_05971_ net139 net1151 _03440_ _03441_ VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__a22o_1
XFILLER_38_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1219 data_array.data0\[5\]\[10\] VGND VGND VPWR VPWR net2870 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_144_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07710_ data_array.data1\[8\]\[24\] net1396 net1302 data_array.data1\[11\]\[24\]
+ _04926_ VGND VGND VPWR VPWR _04927_ sky130_fd_sc_hd__a221o_1
Xfanout1570 net1573 VGND VGND VPWR VPWR net1570 sky130_fd_sc_hd__clkbuf_4
X_08690_ net2528 net764 net487 VGND VGND VPWR VPWR _00449_ sky130_fd_sc_hd__mux2_1
XFILLER_38_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1581 net1582 VGND VGND VPWR VPWR net1581 sky130_fd_sc_hd__clkbuf_4
Xfanout1592 net1594 VGND VGND VPWR VPWR net1592 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_105_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07641_ data_array.data1\[5\]\[18\] net1536 net1440 data_array.data1\[6\]\[18\] VGND
+ VGND VPWR VPWR _04864_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_140_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07572_ _04800_ _04801_ VGND VGND VPWR VPWR _00066_ sky130_fd_sc_hd__or2_2
XFILLER_18_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09311_ net734 net4251 net543 VGND VGND VPWR VPWR _01065_ sky130_fd_sc_hd__mux2_1
X_06523_ tag_array.tag1\[5\]\[5\] net1611 net1515 tag_array.tag1\[6\]\[5\] VGND VGND
+ VPWR VPWR _03848_ sky130_fd_sc_hd__a22o_1
XFILLER_22_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09242_ net713 net3255 net645 VGND VGND VPWR VPWR _00996_ sky130_fd_sc_hd__mux2_1
XFILLER_21_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06454_ tag_array.tag0\[0\]\[24\] net1372 net1278 tag_array.tag0\[3\]\[24\] _03784_
+ VGND VGND VPWR VPWR _03785_ sky130_fd_sc_hd__a221o_1
XFILLER_178_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09173_ net789 net2822 net627 VGND VGND VPWR VPWR _00927_ sky130_fd_sc_hd__mux2_1
X_06385_ tag_array.tag0\[13\]\[18\] net1565 net1469 tag_array.tag0\[14\]\[18\] VGND
+ VGND VPWR VPWR _03722_ sky130_fd_sc_hd__a22o_1
X_08124_ data_array.data1\[8\]\[62\] net1415 net1321 data_array.data1\[11\]\[62\]
+ _05302_ VGND VGND VPWR VPWR _05303_ sky130_fd_sc_hd__a221o_1
XFILLER_175_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08055_ net1216 _05235_ _05239_ net1168 VGND VGND VPWR VPWR _05241_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_116_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07006_ data_array.data0\[8\]\[24\] net1386 net1292 data_array.data0\[11\]\[24\]
+ _04286_ VGND VGND VPWR VPWR _04287_ sky130_fd_sc_hd__a221o_1
XFILLER_150_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_164_3505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2410 data_array.data0\[15\]\[0\] VGND VGND VPWR VPWR net4061 sky130_fd_sc_hd__dlygate4sd3_1
Xinput106 mem_rdata[16] VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_181_3830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2421 tag_array.tag1\[5\]\[23\] VGND VGND VPWR VPWR net4072 sky130_fd_sc_hd__dlygate4sd3_1
Xinput117 mem_rdata[26] VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__clkbuf_1
Xinput128 mem_rdata[36] VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_181_3841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2432 data_array.data1\[12\]\[52\] VGND VGND VPWR VPWR net4083 sky130_fd_sc_hd__dlygate4sd3_1
Xinput139 mem_rdata[46] VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_1
X_08957_ net936 net3323 net431 VGND VGND VPWR VPWR _00713_ sky130_fd_sc_hd__mux2_1
Xhold2443 data_array.data0\[9\]\[31\] VGND VGND VPWR VPWR net4094 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2454 tag_array.tag1\[9\]\[17\] VGND VGND VPWR VPWR net4105 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1720 data_array.data1\[10\]\[63\] VGND VGND VPWR VPWR net3371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2465 tag_array.tag1\[7\]\[23\] VGND VGND VPWR VPWR net4116 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2476 data_array.data1\[14\]\[7\] VGND VGND VPWR VPWR net4127 sky130_fd_sc_hd__dlygate4sd3_1
X_07908_ data_array.data1\[12\]\[42\] net1399 net1305 data_array.data1\[15\]\[42\]
+ _05106_ VGND VGND VPWR VPWR _05107_ sky130_fd_sc_hd__a221o_1
Xhold1731 data_array.data0\[12\]\[55\] VGND VGND VPWR VPWR net3382 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2487 data_array.data0\[6\]\[51\] VGND VGND VPWR VPWR net4138 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1742 data_array.data0\[9\]\[45\] VGND VGND VPWR VPWR net3393 sky130_fd_sc_hd__dlygate4sd3_1
X_08888_ net954 net4147 net437 VGND VGND VPWR VPWR _00645_ sky130_fd_sc_hd__mux2_1
XFILLER_5_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1753 lru_array.lru_mem\[7\] VGND VGND VPWR VPWR net3404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2498 tag_array.tag0\[6\]\[5\] VGND VGND VPWR VPWR net4149 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1764 data_array.data1\[7\]\[45\] VGND VGND VPWR VPWR net3415 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1775 data_array.data1\[3\]\[26\] VGND VGND VPWR VPWR net3426 sky130_fd_sc_hd__dlygate4sd3_1
X_07839_ data_array.data1\[5\]\[36\] net1604 net1508 data_array.data1\[6\]\[36\] VGND
+ VGND VPWR VPWR _05044_ sky130_fd_sc_hd__a22o_1
XFILLER_44_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1786 data_array.data0\[14\]\[2\] VGND VGND VPWR VPWR net3437 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1797 tag_array.tag1\[5\]\[19\] VGND VGND VPWR VPWR net3448 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_71_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10850_ net1085 net4043 net514 VGND VGND VPWR VPWR _02595_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_179_3792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09509_ net794 net2878 net622 VGND VGND VPWR VPWR _01262_ sky130_fd_sc_hd__mux2_1
XFILLER_169_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10781_ net1871 net1104 net502 VGND VGND VPWR VPWR _02526_ sky130_fd_sc_hd__mux2_1
X_12520_ clknet_leaf_32_clk _01214_ VGND VGND VPWR VPWR tag_array.tag1\[11\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_23_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_117_Right_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12451_ clknet_leaf_19_clk _01145_ VGND VGND VPWR VPWR data_array.data1\[9\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11402_ clknet_leaf_140_clk _00212_ VGND VGND VPWR VPWR tag_array.tag1\[7\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12382_ clknet_leaf_230_clk _01076_ VGND VGND VPWR VPWR data_array.data0\[14\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_90 net1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_895 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14121_ clknet_leaf_91_clk _02750_ VGND VGND VPWR VPWR data_array.data0\[1\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_153_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11333_ net960 net2541 net798 VGND VGND VPWR VPWR _03076_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14052_ clknet_leaf_30_clk _02681_ VGND VGND VPWR VPWR data_array.data1\[6\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_11264_ net975 net4415 net673 VGND VGND VPWR VPWR _03007_ sky130_fd_sc_hd__mux2_1
XFILLER_106_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13003_ clknet_leaf_15_clk _01697_ VGND VGND VPWR VPWR data_array.data0\[3\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_10215_ net946 net4197 net355 VGND VGND VPWR VPWR _01962_ sky130_fd_sc_hd__mux2_1
XFILLER_122_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11195_ net995 net4518 net655 VGND VGND VPWR VPWR _02938_ sky130_fd_sc_hd__mux2_1
X_10146_ net962 net4045 net364 VGND VGND VPWR VPWR _01894_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10077_ net716 net3660 net600 VGND VGND VPWR VPWR _01826_ sky130_fd_sc_hd__mux2_1
XFILLER_48_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13905_ clknet_leaf_57_clk _02534_ VGND VGND VPWR VPWR data_array.data1\[4\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_195_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_195_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_48_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13836_ clknet_leaf_69_clk _02465_ VGND VGND VPWR VPWR data_array.data1\[3\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13767_ clknet_leaf_193_clk _02396_ VGND VGND VPWR VPWR data_array.data1\[1\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
X_10979_ net1927 net1084 net336 VGND VGND VPWR VPWR _02723_ sky130_fd_sc_hd__mux2_1
XFILLER_43_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12718_ clknet_leaf_166_clk _01412_ VGND VGND VPWR VPWR tag_array.tag0\[7\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_13698_ clknet_leaf_203_clk _02327_ VGND VGND VPWR VPWR data_array.data1\[15\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1001 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12649_ clknet_leaf_34_clk _01343_ VGND VGND VPWR VPWR data_array.data0\[15\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_154_Left_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06170_ net29 net28 VGND VGND VPWR VPWR _03527_ sky130_fd_sc_hd__nand2b_1
XFILLER_172_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14319_ clknet_leaf_240_clk _02948_ VGND VGND VPWR VPWR data_array.data1\[11\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold305 data_array.data1\[1\]\[45\] VGND VGND VPWR VPWR net1956 sky130_fd_sc_hd__dlygate4sd3_1
Xhold316 data_array.data1\[8\]\[46\] VGND VGND VPWR VPWR net1967 sky130_fd_sc_hd__dlygate4sd3_1
Xhold327 data_array.data0\[8\]\[60\] VGND VGND VPWR VPWR net1978 sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 data_array.data1\[0\]\[12\] VGND VGND VPWR VPWR net1989 sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 data_array.data1\[0\]\[8\] VGND VGND VPWR VPWR net2000 sky130_fd_sc_hd__dlygate4sd3_1
X_09860_ net1028 net4542 net384 VGND VGND VPWR VPWR _01610_ sky130_fd_sc_hd__mux2_1
Xfanout807 _05415_ VGND VGND VPWR VPWR net807 sky130_fd_sc_hd__clkbuf_4
XFILLER_98_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout818 _05359_ VGND VGND VPWR VPWR net818 sky130_fd_sc_hd__clkbuf_2
XFILLER_140_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_74_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout829 net835 VGND VGND VPWR VPWR net829 sky130_fd_sc_hd__buf_12
XFILLER_58_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08811_ net2232 net1003 net445 VGND VGND VPWR VPWR _00569_ sky130_fd_sc_hd__mux2_1
X_09791_ net1046 net4082 net389 VGND VGND VPWR VPWR _01542_ sky130_fd_sc_hd__mux2_1
XFILLER_97_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1005 data_array.data0\[2\]\[44\] VGND VGND VPWR VPWR net2656 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_163_Left_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1016 data_array.data0\[12\]\[34\] VGND VGND VPWR VPWR net2667 sky130_fd_sc_hd__dlygate4sd3_1
X_08742_ net757 net4350 net463 VGND VGND VPWR VPWR _00501_ sky130_fd_sc_hd__mux2_1
Xhold1027 data_array.data0\[7\]\[52\] VGND VGND VPWR VPWR net2678 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05954_ data_array.rdata0\[41\] net847 net1143 VGND VGND VPWR VPWR _03430_ sky130_fd_sc_hd__o21a_1
Xhold1038 tag_array.tag0\[15\]\[12\] VGND VGND VPWR VPWR net2689 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 tag_array.tag1\[12\]\[16\] VGND VGND VPWR VPWR net2700 sky130_fd_sc_hd__dlygate4sd3_1
X_08673_ net730 net4311 net499 VGND VGND VPWR VPWR _00432_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_186_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_186_clk
+ sky130_fd_sc_hd__clkbuf_8
X_05885_ data_array.rdata0\[18\] net847 net1143 VGND VGND VPWR VPWR _03384_ sky130_fd_sc_hd__o21a_1
X_07624_ data_array.data1\[0\]\[16\] net1353 net1259 data_array.data1\[3\]\[16\] _04848_
+ VGND VGND VPWR VPWR _04849_ sky130_fd_sc_hd__a221o_1
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07555_ data_array.data1\[13\]\[10\] net1604 net1508 data_array.data1\[14\]\[10\]
+ VGND VGND VPWR VPWR _04786_ sky130_fd_sc_hd__a22o_1
X_06506_ tag_array.tag1\[9\]\[4\] net1552 net1456 tag_array.tag1\[10\]\[4\] VGND VGND
+ VPWR VPWR _03832_ sky130_fd_sc_hd__a22o_1
XFILLER_22_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07486_ data_array.data1\[8\]\[4\] net1393 net1299 data_array.data1\[11\]\[4\] _04722_
+ VGND VGND VPWR VPWR _04723_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_157_3375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_3386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_172_Left_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09225_ net781 net2974 net645 VGND VGND VPWR VPWR _00979_ sky130_fd_sc_hd__mux2_1
XFILLER_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06437_ net1626 _03763_ _03767_ net1201 VGND VGND VPWR VPWR _03770_ sky130_fd_sc_hd__a22o_1
XFILLER_107_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_118_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09156_ net918 net4509 net574 VGND VGND VPWR VPWR _00910_ sky130_fd_sc_hd__mux2_1
XFILLER_154_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06368_ tag_array.tag0\[12\]\[16\] net1410 net1316 tag_array.tag0\[15\]\[16\] _03706_
+ VGND VGND VPWR VPWR _03707_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_135_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08107_ data_array.data1\[1\]\[60\] net1604 net1508 data_array.data1\[2\]\[60\] VGND
+ VGND VPWR VPWR _05288_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_135_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09087_ net936 net4341 net415 VGND VGND VPWR VPWR _00841_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_110_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_110_clk
+ sky130_fd_sc_hd__clkbuf_8
X_06299_ tag_array.tag0\[5\]\[10\] net1596 net1500 tag_array.tag0\[6\]\[10\] VGND
+ VGND VPWR VPWR _03644_ sky130_fd_sc_hd__a22o_1
XFILLER_174_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08038_ data_array.data1\[0\]\[54\] net1353 net1259 data_array.data1\[3\]\[54\] _05224_
+ VGND VGND VPWR VPWR _05225_ sky130_fd_sc_hd__a221o_1
XFILLER_107_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold850 tag_array.tag1\[10\]\[7\] VGND VGND VPWR VPWR net2501 sky130_fd_sc_hd__dlygate4sd3_1
Xhold861 data_array.data0\[0\]\[26\] VGND VGND VPWR VPWR net2512 sky130_fd_sc_hd__dlygate4sd3_1
Xhold872 data_array.data1\[5\]\[47\] VGND VGND VPWR VPWR net2523 sky130_fd_sc_hd__dlygate4sd3_1
Xhold883 data_array.data0\[13\]\[2\] VGND VGND VPWR VPWR net2534 sky130_fd_sc_hd__dlygate4sd3_1
Xhold894 data_array.data1\[9\]\[63\] VGND VGND VPWR VPWR net2545 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10000_ net1086 net3748 net554 VGND VGND VPWR VPWR _01749_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_181_Left_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09989_ net872 net3482 net376 VGND VGND VPWR VPWR _01738_ sky130_fd_sc_hd__mux2_1
Xhold2240 tag_array.tag0\[3\]\[7\] VGND VGND VPWR VPWR net3891 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2251 data_array.data1\[7\]\[4\] VGND VGND VPWR VPWR net3902 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2262 data_array.data1\[9\]\[35\] VGND VGND VPWR VPWR net3913 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_5_5__f_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_5_5__leaf_clk sky130_fd_sc_hd__clkbuf_16
Xhold2273 data_array.data0\[10\]\[58\] VGND VGND VPWR VPWR net3924 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_92_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2284 data_array.data0\[6\]\[56\] VGND VGND VPWR VPWR net3935 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1550 tag_array.tag1\[9\]\[16\] VGND VGND VPWR VPWR net3201 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2295 data_array.data0\[3\]\[14\] VGND VGND VPWR VPWR net3946 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1561 tag_array.tag0\[3\]\[15\] VGND VGND VPWR VPWR net3212 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1572 data_array.data0\[3\]\[30\] VGND VGND VPWR VPWR net3223 sky130_fd_sc_hd__dlygate4sd3_1
X_11951_ clknet_leaf_268_clk _00759_ VGND VGND VPWR VPWR data_array.data0\[4\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_177_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_177_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold1583 data_array.data0\[15\]\[24\] VGND VGND VPWR VPWR net3234 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_28_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1594 data_array.data1\[12\]\[35\] VGND VGND VPWR VPWR net3245 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_28_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10902_ net878 net2957 net517 VGND VGND VPWR VPWR _02647_ sky130_fd_sc_hd__mux2_1
X_11882_ clknet_leaf_127_clk _00690_ VGND VGND VPWR VPWR data_array.data0\[5\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_10833_ net2315 net898 net502 VGND VGND VPWR VPWR _02578_ sky130_fd_sc_hd__mux2_1
X_13621_ clknet_leaf_23_clk _02250_ VGND VGND VPWR VPWR data_array.data0\[9\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10764_ net918 net4275 net497 VGND VGND VPWR VPWR _02509_ sky130_fd_sc_hd__mux2_1
X_13552_ clknet_leaf_56_clk _02181_ VGND VGND VPWR VPWR data_array.data1\[0\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
X_12503_ clknet_leaf_17_clk _01197_ VGND VGND VPWR VPWR data_array.data1\[9\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_157_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13483_ clknet_leaf_170_clk _02113_ VGND VGND VPWR VPWR tag_array.tag0\[15\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_698 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10695_ net4464 net937 net483 VGND VGND VPWR VPWR _02440_ sky130_fd_sc_hd__mux2_1
XFILLER_139_862 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12434_ clknet_leaf_224_clk _01128_ VGND VGND VPWR VPWR data_array.data0\[14\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_126_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12365_ clknet_leaf_77_clk _00041_ VGND VGND VPWR VPWR data_array.rdata0\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_172_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_101_clk clknet_5_24__leaf_clk VGND VGND VPWR VPWR clknet_leaf_101_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_126_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11316_ net1030 net3836 net805 VGND VGND VPWR VPWR _03059_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14104_ clknet_leaf_222_clk _02733_ VGND VGND VPWR VPWR data_array.data0\[1\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12296_ clknet_leaf_191_clk _01054_ VGND VGND VPWR VPWR tag_array.tag1\[12\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14035_ clknet_leaf_35_clk _02664_ VGND VGND VPWR VPWR data_array.data1\[6\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_11247_ net1041 net3816 net674 VGND VGND VPWR VPWR _02990_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11178_ net1063 net3763 net657 VGND VGND VPWR VPWR _02921_ sky130_fd_sc_hd__mux2_1
XFILLER_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10129_ net1029 net2945 net368 VGND VGND VPWR VPWR _01877_ sky130_fd_sc_hd__mux2_1
XFILLER_94_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_168_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_168_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_91_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_05670_ fsm.tag_out0\[10\] net9 VGND VGND VPWR VPWR _03187_ sky130_fd_sc_hd__and2b_1
XFILLER_51_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13819_ clknet_leaf_4_clk _02448_ VGND VGND VPWR VPWR data_array.data1\[2\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07340_ net1218 _04585_ _04589_ net1170 VGND VGND VPWR VPWR _04591_ sky130_fd_sc_hd__a22o_1
XFILLER_32_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07271_ data_array.data0\[1\]\[48\] net1572 net1476 data_array.data0\[2\]\[48\] VGND
+ VGND VPWR VPWR _04528_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_14_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09010_ net1806 net987 net423 VGND VGND VPWR VPWR _00765_ sky130_fd_sc_hd__mux2_1
X_06222_ tag_array.tag0\[1\]\[3\] net1561 net1465 tag_array.tag0\[2\]\[3\] VGND VGND
+ VPWR VPWR _03574_ sky130_fd_sc_hd__a22o_1
XFILLER_89_1030 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_152_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06153_ net26 net27 VGND VGND VPWR VPWR _03510_ sky130_fd_sc_hd__and2b_1
XFILLER_8_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold102 data_array.data0\[0\]\[15\] VGND VGND VPWR VPWR net1753 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold113 data_array.data0\[2\]\[22\] VGND VGND VPWR VPWR net1764 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold124 data_array.data0\[2\]\[50\] VGND VGND VPWR VPWR net1775 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_567 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold135 data_array.data0\[4\]\[24\] VGND VGND VPWR VPWR net1786 sky130_fd_sc_hd__dlygate4sd3_1
X_06084_ fsm.tag_out0\[24\] net1120 _03505_ VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__a21o_1
Xhold146 data_array.data0\[1\]\[33\] VGND VGND VPWR VPWR net1797 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 tag_array.tag1\[1\]\[19\] VGND VGND VPWR VPWR net1808 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 data_array.data0\[1\]\[13\] VGND VGND VPWR VPWR net1819 sky130_fd_sc_hd__dlygate4sd3_1
X_09912_ net758 net3807 net604 VGND VGND VPWR VPWR _01662_ sky130_fd_sc_hd__mux2_1
Xhold179 data_array.data0\[2\]\[42\] VGND VGND VPWR VPWR net1830 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout604 _05582_ VGND VGND VPWR VPWR net604 sky130_fd_sc_hd__buf_4
Xfanout615 _05571_ VGND VGND VPWR VPWR net615 sky130_fd_sc_hd__buf_4
Xfanout626 _05565_ VGND VGND VPWR VPWR net626 sky130_fd_sc_hd__buf_2
XFILLER_113_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout637 net638 VGND VGND VPWR VPWR net637 sky130_fd_sc_hd__clkbuf_8
X_09843_ net1097 net2583 net382 VGND VGND VPWR VPWR _01593_ sky130_fd_sc_hd__mux2_1
Xfanout648 net651 VGND VGND VPWR VPWR net648 sky130_fd_sc_hd__buf_4
Xfanout659 net660 VGND VGND VPWR VPWR net659 sky130_fd_sc_hd__buf_4
XFILLER_58_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06986_ data_array.data0\[4\]\[22\] net1340 net1246 data_array.data0\[7\]\[22\] _04268_
+ VGND VGND VPWR VPWR _04269_ sky130_fd_sc_hd__a221o_1
X_09774_ net807 _05561_ VGND VGND VPWR VPWR _03125_ sky130_fd_sc_hd__nand2_1
XFILLER_100_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08725_ net2504 net724 net475 VGND VGND VPWR VPWR _00484_ sky130_fd_sc_hd__mux2_1
X_05937_ data_array.rdata1\[35\] net828 net837 VGND VGND VPWR VPWR _03419_ sky130_fd_sc_hd__a21o_1
XFILLER_27_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_159_clk clknet_5_28__leaf_clk VGND VGND VPWR VPWR clknet_leaf_159_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_2_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08656_ net3486 net700 net511 VGND VGND VPWR VPWR _00415_ sky130_fd_sc_hd__mux2_1
X_05868_ data_array.rdata1\[12\] net834 net843 VGND VGND VPWR VPWR _03373_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_159_3415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07607_ data_array.data1\[8\]\[15\] net1394 net1300 data_array.data1\[11\]\[15\]
+ _04832_ VGND VGND VPWR VPWR _04833_ sky130_fd_sc_hd__a221o_1
XFILLER_14_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08587_ net775 net2598 net528 VGND VGND VPWR VPWR _00346_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_176_3740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05799_ _03182_ _03184_ _03200_ _03209_ VGND VGND VPWR VPWR _03316_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_176_3751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07538_ net1168 _04765_ _04769_ net1216 VGND VGND VPWR VPWR _04771_ sky130_fd_sc_hd__a22o_1
XFILLER_23_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07469_ data_array.data1\[1\]\[2\] net1530 net1434 data_array.data1\[2\]\[2\] VGND
+ VGND VPWR VPWR _04708_ sky130_fd_sc_hd__a22o_1
X_09208_ net749 net2726 net630 VGND VGND VPWR VPWR _00962_ sky130_fd_sc_hd__mux2_1
X_10480_ net1026 net4319 net347 VGND VGND VPWR VPWR _02225_ sky130_fd_sc_hd__mux2_1
XFILLER_136_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09139_ net985 net3802 net573 VGND VGND VPWR VPWR _00893_ sky130_fd_sc_hd__mux2_1
X_12150_ clknet_leaf_158_clk _00958_ VGND VGND VPWR VPWR tag_array.tag0\[13\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_108_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11101_ net2333 net857 net330 VGND VGND VPWR VPWR _02844_ sky130_fd_sc_hd__mux2_1
XFILLER_118_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12081_ clknet_leaf_248_clk _00889_ VGND VGND VPWR VPWR data_array.data1\[14\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_123_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold680 tag_array.tag1\[0\]\[18\] VGND VGND VPWR VPWR net2331 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold691 data_array.data1\[9\]\[45\] VGND VGND VPWR VPWR net2342 sky130_fd_sc_hd__dlygate4sd3_1
X_11032_ net2267 net872 net342 VGND VGND VPWR VPWR _02776_ sky130_fd_sc_hd__mux2_1
XFILLER_78_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2070 data_array.data0\[10\]\[26\] VGND VGND VPWR VPWR net3721 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2081 data_array.data1\[14\]\[30\] VGND VGND VPWR VPWR net3732 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2092 data_array.data0\[3\]\[35\] VGND VGND VPWR VPWR net3743 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_94_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12983_ clknet_leaf_159_clk _01677_ VGND VGND VPWR VPWR tag_array.tag0\[4\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_100_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1380 data_array.data1\[13\]\[20\] VGND VGND VPWR VPWR net3031 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1391 data_array.data0\[15\]\[5\] VGND VGND VPWR VPWR net3042 sky130_fd_sc_hd__dlygate4sd3_1
X_11934_ clknet_leaf_16_clk _00742_ VGND VGND VPWR VPWR data_array.data0\[4\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11865_ clknet_leaf_48_clk _00673_ VGND VGND VPWR VPWR data_array.data0\[5\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_13604_ clknet_leaf_54_clk _02233_ VGND VGND VPWR VPWR data_array.data0\[9\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_10816_ net2161 net966 net510 VGND VGND VPWR VPWR _02561_ sky130_fd_sc_hd__mux2_1
X_11796_ clknet_leaf_124_clk _00604_ VGND VGND VPWR VPWR data_array.data0\[8\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
X_13535_ clknet_leaf_257_clk _02164_ VGND VGND VPWR VPWR data_array.data1\[0\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_41_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10747_ net984 net2898 net496 VGND VGND VPWR VPWR _02492_ sky130_fd_sc_hd__mux2_1
XFILLER_174_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10678_ net2111 net1005 net480 VGND VGND VPWR VPWR _02423_ sky130_fd_sc_hd__mux2_1
X_13466_ clknet_leaf_191_clk _02096_ VGND VGND VPWR VPWR tag_array.tag0\[1\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_174_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12417_ clknet_leaf_241_clk _01111_ VGND VGND VPWR VPWR data_array.data0\[14\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_58_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13397_ clknet_leaf_251_clk _02027_ VGND VGND VPWR VPWR data_array.data1\[8\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput207 net207 VGND VGND VPWR VPWR cpu_rdata[48] sky130_fd_sc_hd__clkbuf_4
Xoutput218 net218 VGND VGND VPWR VPWR cpu_rdata[58] sky130_fd_sc_hd__clkbuf_4
XFILLER_182_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12348_ clknet_leaf_68_clk _00023_ VGND VGND VPWR VPWR data_array.rdata0\[30\] sky130_fd_sc_hd__dfxtp_1
Xoutput229 net229 VGND VGND VPWR VPWR cpu_ready sky130_fd_sc_hd__buf_2
XFILLER_114_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12279_ clknet_leaf_33_clk _01037_ VGND VGND VPWR VPWR tag_array.tag1\[13\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14018_ clknet_leaf_201_clk _02647_ VGND VGND VPWR VPWR data_array.data1\[5\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_71_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06840_ data_array.data0\[13\]\[9\] net1580 net1484 data_array.data0\[14\]\[9\] VGND
+ VGND VPWR VPWR _04136_ sky130_fd_sc_hd__a22o_1
XFILLER_96_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_476 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06771_ data_array.data0\[12\]\[3\] net1377 net1283 data_array.data0\[15\]\[3\] _04072_
+ VGND VGND VPWR VPWR _04073_ sky130_fd_sc_hd__a221o_1
X_08510_ _03509_ _03527_ VGND VGND VPWR VPWR _05577_ sky130_fd_sc_hd__nor2_1
X_05722_ net32 fsm.tag_out1\[2\] VGND VGND VPWR VPWR _03239_ sky130_fd_sc_hd__xor2_1
X_09490_ net769 net3879 net624 VGND VGND VPWR VPWR _01243_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08441_ net2205 net888 net687 VGND VGND VPWR VPWR _00276_ sky130_fd_sc_hd__mux2_1
XFILLER_91_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05653_ fsm.tag_out0\[3\] net2 VGND VGND VPWR VPWR _03170_ sky130_fd_sc_hd__and2b_1
XFILLER_23_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08372_ net2457 net982 net686 VGND VGND VPWR VPWR _00253_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_154_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07323_ data_array.data0\[0\]\[53\] net1334 net1240 data_array.data0\[3\]\[53\] _04574_
+ VGND VGND VPWR VPWR _04575_ sky130_fd_sc_hd__a221o_1
XFILLER_20_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_1016 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07254_ data_array.data0\[9\]\[47\] net1577 net1481 data_array.data0\[10\]\[47\]
+ VGND VGND VPWR VPWR _04512_ sky130_fd_sc_hd__a22o_1
XFILLER_164_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06205_ tag_array.tag0\[0\]\[1\] net1401 net1307 tag_array.tag0\[3\]\[1\] _03558_
+ VGND VGND VPWR VPWR _03559_ sky130_fd_sc_hd__a221o_1
X_07185_ net1209 _04443_ _04447_ net1635 VGND VGND VPWR VPWR _04450_ sky130_fd_sc_hd__a22o_1
XFILLER_117_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06136_ data_array.rdata0\[51\] net1134 net1112 data_array.rdata1\[51\] VGND VGND
+ VPWR VPWR net309 sky130_fd_sc_hd__a22o_1
XFILLER_145_695 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06067_ net1163 net16 fsm.tag_out1\[16\] net1133 VGND VGND VPWR VPWR _03497_ sky130_fd_sc_hd__a22o_1
XFILLER_132_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout401 _03124_ VGND VGND VPWR VPWR net401 sky130_fd_sc_hd__buf_4
Xfanout412 net413 VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__buf_4
XFILLER_48_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout423 net425 VGND VGND VPWR VPWR net423 sky130_fd_sc_hd__buf_4
XFILLER_120_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout434 net441 VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__clkbuf_8
XFILLER_87_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout445 net449 VGND VGND VPWR VPWR net445 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout456 net459 VGND VGND VPWR VPWR net456 sky130_fd_sc_hd__clkbuf_4
X_09826_ net905 net4130 net386 VGND VGND VPWR VPWR _01577_ sky130_fd_sc_hd__mux2_1
XFILLER_59_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout467 net468 VGND VGND VPWR VPWR net467 sky130_fd_sc_hd__clkbuf_8
XFILLER_100_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout478 net480 VGND VGND VPWR VPWR net478 sky130_fd_sc_hd__clkbuf_8
Xfanout489 _05602_ VGND VGND VPWR VPWR net489 sky130_fd_sc_hd__clkbuf_4
XFILLER_87_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09757_ net1941 net760 net672 VGND VGND VPWR VPWR _01509_ sky130_fd_sc_hd__mux2_1
X_06969_ data_array.data0\[8\]\[21\] net1365 net1271 data_array.data0\[11\]\[21\]
+ _04252_ VGND VGND VPWR VPWR _04253_ sky130_fd_sc_hd__a221o_1
XFILLER_27_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08708_ net1888 net791 net471 VGND VGND VPWR VPWR _00467_ sky130_fd_sc_hd__mux2_1
X_09688_ net736 net3553 net605 VGND VGND VPWR VPWR _01440_ sky130_fd_sc_hd__mux2_1
XFILLER_15_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08639_ net2377 net766 net513 VGND VGND VPWR VPWR _00398_ sky130_fd_sc_hd__mux2_1
XFILLER_81_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_855 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11650_ clknet_leaf_140_clk _00458_ VGND VGND VPWR VPWR tag_array.tag1\[2\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10601_ net1787 net1056 net469 VGND VGND VPWR VPWR _02346_ sky130_fd_sc_hd__mux2_1
XFILLER_70_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11581_ clknet_leaf_194_clk _00389_ VGND VGND VPWR VPWR tag_array.tag1\[5\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_156_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_915 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10532_ net1078 net4376 net455 VGND VGND VPWR VPWR _02277_ sky130_fd_sc_hd__mux2_1
X_13320_ clknet_leaf_54_clk _01950_ VGND VGND VPWR VPWR data_array.data0\[10\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10463_ net1093 net3794 net349 VGND VGND VPWR VPWR _02208_ sky130_fd_sc_hd__mux2_1
X_13251_ clknet_leaf_96_clk _01881_ VGND VGND VPWR VPWR data_array.data0\[11\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_170_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12202_ clknet_leaf_148_clk _00155_ VGND VGND VPWR VPWR fsm.tag_out0\[9\] sky130_fd_sc_hd__dfxtp_2
X_13182_ clknet_leaf_67_clk _00074_ VGND VGND VPWR VPWR data_array.rdata1\[19\] sky130_fd_sc_hd__dfxtp_1
X_10394_ net2000 net1078 net663 VGND VGND VPWR VPWR _02140_ sky130_fd_sc_hd__mux2_1
X_12133_ clknet_leaf_162_clk _00941_ VGND VGND VPWR VPWR tag_array.tag0\[12\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_53_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12064_ clknet_leaf_119_clk _00872_ VGND VGND VPWR VPWR data_array.data1\[14\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_89_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11015_ net2276 net940 net343 VGND VGND VPWR VPWR _02759_ sky130_fd_sc_hd__mux2_1
XFILLER_77_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout990 _05480_ VGND VGND VPWR VPWR net990 sky130_fd_sc_hd__clkbuf_2
XFILLER_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12966_ clknet_leaf_181_clk _01660_ VGND VGND VPWR VPWR tag_array.tag0\[4\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_16_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11917_ clknet_leaf_14_clk _00725_ VGND VGND VPWR VPWR data_array.data0\[5\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12897_ clknet_leaf_261_clk _01591_ VGND VGND VPWR VPWR data_array.data0\[13\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_61_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11848_ clknet_leaf_25_clk _00656_ VGND VGND VPWR VPWR data_array.data0\[7\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11779_ clknet_leaf_27_clk _00587_ VGND VGND VPWR VPWR data_array.data0\[8\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13518_ clknet_leaf_64_clk _02147_ VGND VGND VPWR VPWR data_array.data1\[0\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_118_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14498_ clknet_leaf_179_clk _03120_ VGND VGND VPWR VPWR lru_array.lru_mem\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_174_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload11 clknet_5_25__leaf_clk VGND VGND VPWR VPWR clkload11/X sky130_fd_sc_hd__clkbuf_8
Xclkload22 clknet_leaf_261_clk VGND VGND VPWR VPWR clkload22/X sky130_fd_sc_hd__clkbuf_8
X_13449_ clknet_leaf_142_clk _02079_ VGND VGND VPWR VPWR tag_array.tag0\[1\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_173_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload33 clknet_leaf_13_clk VGND VGND VPWR VPWR clkload33/Y sky130_fd_sc_hd__inv_6
Xclkload44 clknet_leaf_244_clk VGND VGND VPWR VPWR clkload44/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload55 clknet_leaf_253_clk VGND VGND VPWR VPWR clkload55/Y sky130_fd_sc_hd__bufinv_16
XFILLER_127_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload66 clknet_leaf_30_clk VGND VGND VPWR VPWR clkload66/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload77 clknet_leaf_49_clk VGND VGND VPWR VPWR clkload77/X sky130_fd_sc_hd__clkbuf_8
Xclkload88 clknet_leaf_53_clk VGND VGND VPWR VPWR clkload88/X sky130_fd_sc_hd__clkbuf_8
XFILLER_170_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload99 clknet_leaf_69_clk VGND VGND VPWR VPWR clkload99/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_126_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08990_ net2211 net1065 net423 VGND VGND VPWR VPWR _00745_ sky130_fd_sc_hd__mux2_1
XFILLER_173_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07941_ data_array.data1\[8\]\[45\] net1350 net1256 data_array.data1\[11\]\[45\]
+ _05136_ VGND VGND VPWR VPWR _05137_ sky130_fd_sc_hd__a221o_1
Xhold2806 data_array.data0\[15\]\[3\] VGND VGND VPWR VPWR net4457 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2817 tag_array.dirty0\[1\] VGND VGND VPWR VPWR net4468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2828 tag_array.tag1\[7\]\[16\] VGND VGND VPWR VPWR net4479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2839 data_array.data1\[7\]\[28\] VGND VGND VPWR VPWR net4490 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_147_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07872_ data_array.data1\[1\]\[39\] net1538 net1442 data_array.data1\[2\]\[39\] VGND
+ VGND VPWR VPWR _05074_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_147_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09611_ net905 net3782 net394 VGND VGND VPWR VPWR _01363_ sky130_fd_sc_hd__mux2_1
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06823_ net1231 _04115_ _04119_ net1183 VGND VGND VPWR VPWR _04121_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_108_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06754_ data_array.data0\[5\]\[1\] net1520 net1424 data_array.data0\[6\]\[1\] VGND
+ VGND VPWR VPWR _04058_ sky130_fd_sc_hd__a22o_1
X_09542_ net758 net2981 net619 VGND VGND VPWR VPWR _01295_ sky130_fd_sc_hd__mux2_1
X_05705_ _03220_ _03221_ _03180_ _03210_ VGND VGND VPWR VPWR _03222_ sky130_fd_sc_hd__a211o_1
X_09473_ net734 net4386 net654 VGND VGND VPWR VPWR _01226_ sky130_fd_sc_hd__mux2_1
X_06685_ tag_array.tag1\[0\]\[20\] net1349 net1255 tag_array.tag1\[3\]\[20\] _03994_
+ VGND VGND VPWR VPWR _03995_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_90_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_90_clk sky130_fd_sc_hd__clkbuf_8
X_08424_ net144 net79 net1642 VGND VGND VPWR VPWR _05519_ sky130_fd_sc_hd__mux2_1
X_05636_ net1649 net1160 net33 VGND VGND VPWR VPWR _03153_ sky130_fd_sc_hd__and3_4
XFILLER_180_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08355_ net118 net53 net1643 VGND VGND VPWR VPWR _05473_ sky130_fd_sc_hd__mux2_1
X_07306_ net1188 _04553_ _04557_ net1615 VGND VGND VPWR VPWR _04560_ sky130_fd_sc_hd__a22o_1
Xclkload5 clknet_5_10__leaf_clk VGND VGND VPWR VPWR clkload5/X sky130_fd_sc_hd__clkbuf_8
X_08286_ net143 net78 net1641 VGND VGND VPWR VPWR _05427_ sky130_fd_sc_hd__mux2_1
XFILLER_137_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07237_ data_array.data0\[8\]\[45\] net1344 net1250 data_array.data0\[11\]\[45\]
+ _04496_ VGND VGND VPWR VPWR _04497_ sky130_fd_sc_hd__a221o_1
XFILLER_166_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07168_ data_array.data0\[1\]\[39\] net1538 net1442 data_array.data0\[2\]\[39\] VGND
+ VGND VPWR VPWR _04434_ sky130_fd_sc_hd__a22o_1
XFILLER_105_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_5_30__f_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_5_30__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_06119_ data_array.rdata0\[34\] net1138 net1113 data_array.rdata1\[34\] VGND VGND
+ VPWR VPWR net290 sky130_fd_sc_hd__a22o_1
X_07099_ _04370_ _04371_ VGND VGND VPWR VPWR _00025_ sky130_fd_sc_hd__or2_1
XFILLER_59_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_3569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1207 net1208 VGND VGND VPWR VPWR net1207 sky130_fd_sc_hd__buf_4
XFILLER_121_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1218 net1220 VGND VGND VPWR VPWR net1218 sky130_fd_sc_hd__buf_4
Xfanout1229 net1230 VGND VGND VPWR VPWR net1229 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_184_3894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09809_ net973 net2667 net386 VGND VGND VPWR VPWR _01560_ sky130_fd_sc_hd__mux2_1
XFILLER_75_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12820_ clknet_leaf_134_clk _01514_ VGND VGND VPWR VPWR tag_array.tag1\[0\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_55_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12751_ clknet_leaf_106_clk _01445_ VGND VGND VPWR VPWR tag_array.tag0\[5\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_81_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_81_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_15_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11702_ clknet_leaf_187_clk _00510_ VGND VGND VPWR VPWR tag_array.tag1\[15\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_131_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12682_ clknet_leaf_106_clk _01376_ VGND VGND VPWR VPWR tag_array.tag0\[8\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14421_ clknet_leaf_198_clk _03044_ VGND VGND VPWR VPWR data_array.data1\[7\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_46_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ clknet_leaf_188_clk _00441_ VGND VGND VPWR VPWR tag_array.tag1\[3\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_1060 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14352_ clknet_leaf_251_clk _02975_ VGND VGND VPWR VPWR data_array.data1\[10\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11564_ clknet_leaf_129_clk _00372_ VGND VGND VPWR VPWR tag_array.tag1\[5\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_763 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13303_ clknet_leaf_94_clk _01933_ VGND VGND VPWR VPWR data_array.data0\[10\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_156_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10515_ net885 net4277 net344 VGND VGND VPWR VPWR _02260_ sky130_fd_sc_hd__mux2_1
XFILLER_128_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11495_ clknet_leaf_172_clk _00304_ VGND VGND VPWR VPWR tag_array.valid1\[9\] sky130_fd_sc_hd__dfxtp_1
X_14283_ clknet_leaf_19_clk _02912_ VGND VGND VPWR VPWR data_array.data1\[11\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10446_ net2101 net870 net671 VGND VGND VPWR VPWR _02192_ sky130_fd_sc_hd__mux2_1
X_13234_ clknet_leaf_94_clk _01864_ VGND VGND VPWR VPWR data_array.data0\[11\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_90_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13165_ clknet_leaf_252_clk _00086_ VGND VGND VPWR VPWR data_array.rdata1\[2\] sky130_fd_sc_hd__dfxtp_1
X_10377_ net824 net1645 VGND VGND VPWR VPWR _03130_ sky130_fd_sc_hd__and2b_2
XFILLER_124_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12116_ clknet_leaf_121_clk _00924_ VGND VGND VPWR VPWR data_array.data1\[14\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
X_13096_ clknet_leaf_77_clk _01790_ VGND VGND VPWR VPWR data_array.data1\[13\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_123_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12047_ clknet_leaf_237_clk _00855_ VGND VGND VPWR VPWR data_array.data0\[6\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_66_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13998_ clknet_leaf_74_clk _02627_ VGND VGND VPWR VPWR data_array.data1\[5\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_142_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12949_ clknet_leaf_3_clk _01643_ VGND VGND VPWR VPWR data_array.data0\[13\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_66_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_72_clk clknet_5_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_72_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_103_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06470_ net1629 _03793_ _03797_ net1203 VGND VGND VPWR VPWR _03800_ sky130_fd_sc_hd__a22o_1
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08140_ data_array.data1\[1\]\[63\] net1553 net1457 data_array.data1\[2\]\[63\] VGND
+ VGND VPWR VPWR _05318_ sky130_fd_sc_hd__a22o_1
XFILLER_14_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload100 clknet_leaf_70_clk VGND VGND VPWR VPWR clkload100/Y sky130_fd_sc_hd__clkinv_2
X_08071_ data_array.data1\[0\]\[57\] net1338 net1244 data_array.data1\[3\]\[57\] _05254_
+ VGND VGND VPWR VPWR _05255_ sky130_fd_sc_hd__a221o_1
Xclkload111 clknet_leaf_94_clk VGND VGND VPWR VPWR clkload111/X sky130_fd_sc_hd__clkbuf_4
Xclkload122 clknet_leaf_89_clk VGND VGND VPWR VPWR clkload122/Y sky130_fd_sc_hd__inv_6
X_07022_ _04300_ _04301_ VGND VGND VPWR VPWR _00017_ sky130_fd_sc_hd__or2_1
Xclkload133 clknet_leaf_215_clk VGND VGND VPWR VPWR clkload133/Y sky130_fd_sc_hd__bufinv_16
XFILLER_174_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload144 clknet_leaf_209_clk VGND VGND VPWR VPWR clkload144/Y sky130_fd_sc_hd__clkinv_8
Xclkload155 clknet_leaf_232_clk VGND VGND VPWR VPWR clkload155/Y sky130_fd_sc_hd__inv_6
Xclkload166 clknet_leaf_204_clk VGND VGND VPWR VPWR clkload166/X sky130_fd_sc_hd__clkbuf_8
XFILLER_161_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload177 clknet_leaf_177_clk VGND VGND VPWR VPWR clkload177/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_149_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload188 clknet_leaf_189_clk VGND VGND VPWR VPWR clkload188/Y sky130_fd_sc_hd__clkinv_2
Xclkload199 clknet_leaf_160_clk VGND VGND VPWR VPWR clkload199/Y sky130_fd_sc_hd__clkinv_2
XFILLER_142_440 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2603 data_array.data1\[10\]\[18\] VGND VGND VPWR VPWR net4254 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08973_ net872 net2972 net430 VGND VGND VPWR VPWR _00729_ sky130_fd_sc_hd__mux2_1
Xhold2614 tag_array.tag0\[7\]\[2\] VGND VGND VPWR VPWR net4265 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_114_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2625 data_array.data1\[12\]\[47\] VGND VGND VPWR VPWR net4276 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2636 data_array.data0\[9\]\[27\] VGND VGND VPWR VPWR net4287 sky130_fd_sc_hd__dlygate4sd3_1
X_07924_ _05120_ _05121_ VGND VGND VPWR VPWR _00101_ sky130_fd_sc_hd__or2_1
Xhold1902 tag_array.tag0\[5\]\[14\] VGND VGND VPWR VPWR net3553 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2647 tag_array.tag0\[4\]\[2\] VGND VGND VPWR VPWR net4298 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2658 data_array.data1\[10\]\[36\] VGND VGND VPWR VPWR net4309 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1913 tag_array.tag0\[12\]\[2\] VGND VGND VPWR VPWR net3564 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1924 data_array.data1\[9\]\[21\] VGND VGND VPWR VPWR net3575 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2669 data_array.data0\[14\]\[3\] VGND VGND VPWR VPWR net4320 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1935 data_array.data1\[5\]\[33\] VGND VGND VPWR VPWR net3586 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_162_3477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07855_ data_array.data1\[4\]\[37\] net1353 net1259 data_array.data1\[7\]\[37\] _05058_
+ VGND VGND VPWR VPWR _05059_ sky130_fd_sc_hd__a221o_1
Xhold1946 data_array.data1\[3\]\[5\] VGND VGND VPWR VPWR net3597 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1957 data_array.data0\[13\]\[36\] VGND VGND VPWR VPWR net3608 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_68_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1968 tag_array.tag0\[11\]\[8\] VGND VGND VPWR VPWR net3619 sky130_fd_sc_hd__dlygate4sd3_1
X_06806_ data_array.data0\[0\]\[6\] net1329 net1235 data_array.data0\[3\]\[6\] _04104_
+ VGND VGND VPWR VPWR _04105_ sky130_fd_sc_hd__a221o_1
Xhold1979 tag_array.tag0\[9\]\[7\] VGND VGND VPWR VPWR net3630 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_123_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07786_ data_array.data1\[9\]\[31\] net1577 net1481 data_array.data1\[10\]\[31\]
+ VGND VGND VPWR VPWR _04996_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_123_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09525_ net726 net3269 net623 VGND VGND VPWR VPWR _01278_ sky130_fd_sc_hd__mux2_1
X_06737_ data_array.data0\[13\]\[0\] net1557 net1461 data_array.data0\[14\]\[0\] VGND
+ VGND VPWR VPWR _04042_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_63_clk clknet_5_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_63_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_25_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06668_ net1200 _03973_ _03977_ net1626 VGND VGND VPWR VPWR _03980_ sky130_fd_sc_hd__a22o_1
X_09456_ net820 net3256 _05566_ VGND VGND VPWR VPWR _01209_ sky130_fd_sc_hd__mux2_1
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08407_ net1129 _05507_ VGND VGND VPWR VPWR _05508_ sky130_fd_sc_hd__and2_1
XFILLER_52_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05619_ fsm.tag_out1\[15\] VGND VGND VPWR VPWR _03141_ sky130_fd_sc_hd__inv_2
XFILLER_12_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09387_ net819 net2221 _05575_ VGND VGND VPWR VPWR _01140_ sky130_fd_sc_hd__mux2_1
X_06599_ tag_array.tag1\[8\]\[12\] net1401 net1307 tag_array.tag1\[11\]\[12\] _03916_
+ VGND VGND VPWR VPWR _03917_ sky130_fd_sc_hd__a221o_1
XFILLER_177_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Left_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08338_ net1125 _05461_ VGND VGND VPWR VPWR _05462_ sky130_fd_sc_hd__and2_1
XFILLER_138_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08269_ fsm.state\[2\] net1644 net840 _05355_ VGND VGND VPWR VPWR _05414_ sky130_fd_sc_hd__a31oi_2
XFILLER_126_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_169_3609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10300_ net2030 net963 net637 VGND VGND VPWR VPWR _02047_ sky130_fd_sc_hd__mux2_1
XFILLER_153_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11280_ net911 net3960 net674 VGND VGND VPWR VPWR _03023_ sky130_fd_sc_hd__mux2_1
XFILLER_152_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10231_ net880 net3469 net357 VGND VGND VPWR VPWR _01978_ sky130_fd_sc_hd__mux2_1
XFILLER_106_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_952 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10162_ net896 net3983 net362 VGND VGND VPWR VPWR _01910_ sky130_fd_sc_hd__mux2_1
XFILLER_117_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1004 net1005 VGND VGND VPWR VPWR net1004 sky130_fd_sc_hd__clkbuf_2
Xfanout1015 _05468_ VGND VGND VPWR VPWR net1015 sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_EDGE_ROW_58_Left_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1026 net1027 VGND VGND VPWR VPWR net1026 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1037 _05456_ VGND VGND VPWR VPWR net1037 sky130_fd_sc_hd__buf_1
X_10093_ net2005 net751 net643 VGND VGND VPWR VPWR _01842_ sky130_fd_sc_hd__mux2_1
Xfanout1048 net1049 VGND VGND VPWR VPWR net1048 sky130_fd_sc_hd__clkbuf_2
Xfanout1059 _05446_ VGND VGND VPWR VPWR net1059 sky130_fd_sc_hd__buf_1
XFILLER_48_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13921_ clknet_leaf_267_clk _02550_ VGND VGND VPWR VPWR data_array.data1\[4\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13852_ clknet_leaf_123_clk _02481_ VGND VGND VPWR VPWR data_array.data1\[3\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12803_ clknet_leaf_102_clk _01497_ VGND VGND VPWR VPWR tag_array.tag1\[10\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13783_ clknet_leaf_64_clk _02412_ VGND VGND VPWR VPWR data_array.data1\[2\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_10995_ net1938 net1020 net337 VGND VGND VPWR VPWR _02739_ sky130_fd_sc_hd__mux2_1
XFILLER_90_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_54_clk clknet_5_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_54_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_37_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12734_ clknet_leaf_168_clk _01428_ VGND VGND VPWR VPWR tag_array.tag0\[5\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_44_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_994 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_67_Left_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12665_ clknet_leaf_38_clk _01359_ VGND VGND VPWR VPWR data_array.data0\[15\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
X_14404_ clknet_leaf_251_clk _03027_ VGND VGND VPWR VPWR data_array.data1\[10\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_61_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11616_ clknet_leaf_132_clk _00424_ VGND VGND VPWR VPWR tag_array.tag1\[3\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_61_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12596_ clknet_leaf_177_clk _01290_ VGND VGND VPWR VPWR tag_array.tag0\[0\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14335_ clknet_leaf_20_clk _02964_ VGND VGND VPWR VPWR data_array.data1\[11\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
X_11547_ clknet_leaf_132_clk _00355_ VGND VGND VPWR VPWR tag_array.tag1\[6\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold509 tag_array.tag1\[1\]\[3\] VGND VGND VPWR VPWR net2160 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_183_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14266_ clknet_leaf_245_clk _02895_ VGND VGND VPWR VPWR data_array.data1\[12\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
X_11478_ clknet_leaf_151_clk _00181_ VGND VGND VPWR VPWR fsm.valid0 sky130_fd_sc_hd__dfxtp_1
X_13217_ clknet_leaf_214_clk _00113_ VGND VGND VPWR VPWR data_array.rdata1\[54\] sky130_fd_sc_hd__dfxtp_1
X_10429_ net1972 net937 net667 VGND VGND VPWR VPWR _02175_ sky130_fd_sc_hd__mux2_1
X_14197_ clknet_leaf_20_clk _02826_ VGND VGND VPWR VPWR data_array.data0\[2\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_76_Left_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13148_ clknet_leaf_105_clk _01842_ VGND VGND VPWR VPWR tag_array.tag1\[8\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_98_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05970_ data_array.rdata1\[46\] net829 net838 VGND VGND VPWR VPWR _03441_ sky130_fd_sc_hd__a21o_1
X_13079_ clknet_leaf_67_clk _01773_ VGND VGND VPWR VPWR data_array.data1\[13\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_25_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1209 data_array.data0\[2\]\[52\] VGND VGND VPWR VPWR net2860 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_144_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1560 net1566 VGND VGND VPWR VPWR net1560 sky130_fd_sc_hd__buf_2
XFILLER_78_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1571 net1573 VGND VGND VPWR VPWR net1571 sky130_fd_sc_hd__clkbuf_2
Xfanout1582 net1591 VGND VGND VPWR VPWR net1582 sky130_fd_sc_hd__clkbuf_4
XFILLER_66_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1593 net1594 VGND VGND VPWR VPWR net1593 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_105_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07640_ data_array.data1\[8\]\[18\] net1345 net1251 data_array.data1\[11\]\[18\]
+ _04862_ VGND VGND VPWR VPWR _04863_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_140_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07571_ net1234 _04795_ _04799_ net1177 VGND VGND VPWR VPWR _04801_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_45_clk clknet_5_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_45_clk sky130_fd_sc_hd__clkbuf_8
X_09310_ net741 net3370 net552 VGND VGND VPWR VPWR _01064_ sky130_fd_sc_hd__mux2_1
X_06522_ tag_array.tag1\[12\]\[5\] net1420 net1326 tag_array.tag1\[15\]\[5\] _03846_
+ VGND VGND VPWR VPWR _03847_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_85_Left_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06453_ tag_array.tag0\[1\]\[24\] net1562 net1466 tag_array.tag0\[2\]\[24\] VGND
+ VGND VPWR VPWR _03784_ sky130_fd_sc_hd__a22o_1
X_09241_ net717 net3621 net646 VGND VGND VPWR VPWR _00995_ sky130_fd_sc_hd__mux2_1
X_09172_ net793 net3581 net628 VGND VGND VPWR VPWR _00926_ sky130_fd_sc_hd__mux2_1
X_06384_ _03720_ _03721_ VGND VGND VPWR VPWR _00139_ sky130_fd_sc_hd__or2_1
XFILLER_119_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08123_ data_array.data1\[9\]\[62\] net1605 net1509 data_array.data1\[10\]\[62\]
+ VGND VGND VPWR VPWR _05302_ sky130_fd_sc_hd__a22o_1
XFILLER_31_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08054_ net1194 _05233_ _05237_ net1620 VGND VGND VPWR VPWR _05240_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_116_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07005_ data_array.data0\[9\]\[24\] net1577 net1481 data_array.data0\[10\]\[24\]
+ VGND VGND VPWR VPWR _04286_ sky130_fd_sc_hd__a22o_1
XFILLER_162_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_164_3506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_164_3517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2400 data_array.data0\[9\]\[14\] VGND VGND VPWR VPWR net4051 sky130_fd_sc_hd__dlygate4sd3_1
Xinput107 mem_rdata[17] VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_1
Xhold2411 data_array.data0\[3\]\[4\] VGND VGND VPWR VPWR net4062 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_181_3831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput118 mem_rdata[27] VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_1
Xhold2422 data_array.data1\[11\]\[45\] VGND VGND VPWR VPWR net4073 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08956_ net940 net3151 net432 VGND VGND VPWR VPWR _00712_ sky130_fd_sc_hd__mux2_1
XFILLER_131_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_181_3842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2433 data_array.data1\[14\]\[42\] VGND VGND VPWR VPWR net4084 sky130_fd_sc_hd__dlygate4sd3_1
Xinput129 mem_rdata[37] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2444 data_array.data0\[5\]\[41\] VGND VGND VPWR VPWR net4095 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1710 data_array.data1\[7\]\[27\] VGND VGND VPWR VPWR net3361 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2455 tag_array.tag1\[14\]\[1\] VGND VGND VPWR VPWR net4106 sky130_fd_sc_hd__dlygate4sd3_1
X_07907_ data_array.data1\[13\]\[42\] net1589 net1493 data_array.data1\[14\]\[42\]
+ VGND VGND VPWR VPWR _05106_ sky130_fd_sc_hd__a22o_1
Xhold2466 tag_array.tag1\[11\]\[6\] VGND VGND VPWR VPWR net4117 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1721 data_array.data1\[15\]\[29\] VGND VGND VPWR VPWR net3372 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2477 data_array.data0\[11\]\[5\] VGND VGND VPWR VPWR net4128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1732 data_array.data1\[7\]\[35\] VGND VGND VPWR VPWR net3383 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1743 tag_array.tag1\[6\]\[14\] VGND VGND VPWR VPWR net3394 sky130_fd_sc_hd__dlygate4sd3_1
X_08887_ net956 net4339 net438 VGND VGND VPWR VPWR _00644_ sky130_fd_sc_hd__mux2_1
Xhold2488 data_array.data0\[7\]\[63\] VGND VGND VPWR VPWR net4139 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2499 data_array.data0\[9\]\[57\] VGND VGND VPWR VPWR net4150 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1754 tag_array.tag1\[4\]\[12\] VGND VGND VPWR VPWR net3405 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1765 data_array.data1\[7\]\[56\] VGND VGND VPWR VPWR net3416 sky130_fd_sc_hd__dlygate4sd3_1
X_07838_ data_array.data1\[8\]\[36\] net1416 net1322 data_array.data1\[11\]\[36\]
+ _05042_ VGND VGND VPWR VPWR _05043_ sky130_fd_sc_hd__a221o_1
XFILLER_99_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1776 data_array.data1\[14\]\[24\] VGND VGND VPWR VPWR net3427 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1787 data_array.data1\[6\]\[60\] VGND VGND VPWR VPWR net3438 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1798 tag_array.dirty1\[3\] VGND VGND VPWR VPWR net3449 sky130_fd_sc_hd__dlygate4sd3_1
X_07769_ net1224 _04975_ _04979_ net1176 VGND VGND VPWR VPWR _04981_ sky130_fd_sc_hd__a22o_1
XFILLER_60_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_36_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_36_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_53_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09508_ net697 net3283 net624 VGND VGND VPWR VPWR _01261_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_179_3793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10780_ net1936 net1110 net506 VGND VGND VPWR VPWR _02525_ sky130_fd_sc_hd__mux2_1
XFILLER_25_696 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09439_ net911 net4190 net579 VGND VGND VPWR VPWR _01192_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12450_ clknet_leaf_251_clk _01144_ VGND VGND VPWR VPWR data_array.data1\[9\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11401_ clknet_leaf_99_clk _00211_ VGND VGND VPWR VPWR tag_array.tag1\[7\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_12381_ clknet_leaf_211_clk _00059_ VGND VGND VPWR VPWR data_array.rdata0\[63\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_80 net433 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_91 net1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14120_ clknet_leaf_258_clk _02749_ VGND VGND VPWR VPWR data_array.data0\[1\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
X_11332_ net966 net4089 net804 VGND VGND VPWR VPWR _03075_ sky130_fd_sc_hd__mux2_1
XFILLER_67_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14051_ clknet_leaf_220_clk _02680_ VGND VGND VPWR VPWR data_array.data1\[6\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_708 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11263_ net979 net4575 net681 VGND VGND VPWR VPWR _03006_ sky130_fd_sc_hd__mux2_1
XFILLER_180_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13002_ clknet_leaf_250_clk _01696_ VGND VGND VPWR VPWR data_array.data0\[3\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10214_ net949 net2594 net360 VGND VGND VPWR VPWR _01961_ sky130_fd_sc_hd__mux2_1
X_11194_ net997 net4454 net650 VGND VGND VPWR VPWR _02937_ sky130_fd_sc_hd__mux2_1
XFILLER_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10145_ net965 net2872 net368 VGND VGND VPWR VPWR _01893_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10076_ net720 net2963 net601 VGND VGND VPWR VPWR _01825_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_85_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13904_ clknet_leaf_28_clk _02533_ VGND VGND VPWR VPWR data_array.data1\[4\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13835_ clknet_leaf_36_clk _02464_ VGND VGND VPWR VPWR data_array.data1\[3\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_27_clk clknet_5_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_63_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13766_ clknet_leaf_120_clk _02395_ VGND VGND VPWR VPWR data_array.data1\[1\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10978_ net2169 net1088 net338 VGND VGND VPWR VPWR _02722_ sky130_fd_sc_hd__mux2_1
XFILLER_15_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12717_ clknet_leaf_107_clk _01411_ VGND VGND VPWR VPWR tag_array.tag0\[7\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13697_ clknet_leaf_239_clk _02326_ VGND VGND VPWR VPWR data_array.data1\[15\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_148_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12648_ clknet_leaf_71_clk _01342_ VGND VGND VPWR VPWR data_array.data0\[15\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12579_ clknet_leaf_161_clk _01273_ VGND VGND VPWR VPWR tag_array.tag0\[10\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14318_ clknet_leaf_77_clk _02947_ VGND VGND VPWR VPWR data_array.data1\[11\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold306 data_array.data1\[1\]\[8\] VGND VGND VPWR VPWR net1957 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold317 data_array.data1\[0\]\[29\] VGND VGND VPWR VPWR net1968 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold328 data_array.data1\[4\]\[7\] VGND VGND VPWR VPWR net1979 sky130_fd_sc_hd__dlygate4sd3_1
Xhold339 data_array.data0\[4\]\[60\] VGND VGND VPWR VPWR net1990 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_78_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14249_ clknet_leaf_75_clk _02878_ VGND VGND VPWR VPWR data_array.data1\[12\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_125_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout808 _05364_ VGND VGND VPWR VPWR net808 sky130_fd_sc_hd__clkbuf_4
Xfanout819 _05356_ VGND VGND VPWR VPWR net819 sky130_fd_sc_hd__clkbuf_2
X_08810_ net2916 net1007 net442 VGND VGND VPWR VPWR _00568_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_74_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09790_ net1048 net2378 net391 VGND VGND VPWR VPWR _01541_ sky130_fd_sc_hd__mux2_1
XFILLER_86_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1006 data_array.data0\[10\]\[24\] VGND VGND VPWR VPWR net2657 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1017 tag_array.tag0\[13\]\[23\] VGND VGND VPWR VPWR net2668 sky130_fd_sc_hd__dlygate4sd3_1
X_08741_ net760 net3691 net464 VGND VGND VPWR VPWR _00500_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_183_Right_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05953_ net133 net1157 _03428_ _03429_ VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__a22o_1
Xhold1028 data_array.data0\[14\]\[52\] VGND VGND VPWR VPWR net2679 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1039 data_array.data1\[14\]\[4\] VGND VGND VPWR VPWR net2690 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1390 net1392 VGND VGND VPWR VPWR net1390 sky130_fd_sc_hd__clkbuf_2
X_05884_ net107 net1150 _03382_ _03383_ VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__a22o_1
X_08672_ net735 net4208 net494 VGND VGND VPWR VPWR _00431_ sky130_fd_sc_hd__mux2_1
XFILLER_26_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07623_ data_array.data1\[1\]\[16\] net1544 net1448 data_array.data1\[2\]\[16\] VGND
+ VGND VPWR VPWR _04848_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_18_clk clknet_5_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_41_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07554_ data_array.data1\[4\]\[10\] net1414 net1320 data_array.data1\[7\]\[10\] _04784_
+ VGND VGND VPWR VPWR _04785_ sky130_fd_sc_hd__a221o_1
XFILLER_81_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06505_ _03830_ _03831_ VGND VGND VPWR VPWR _00174_ sky130_fd_sc_hd__or2_1
X_07485_ data_array.data1\[9\]\[4\] net1583 net1487 data_array.data1\[10\]\[4\] VGND
+ VGND VPWR VPWR _04722_ sky130_fd_sc_hd__a22o_1
XFILLER_34_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_3376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_3387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_1036 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09224_ net785 net2417 net645 VGND VGND VPWR VPWR _00978_ sky130_fd_sc_hd__mux2_1
X_06436_ tag_array.tag0\[0\]\[22\] net1375 net1281 tag_array.tag0\[3\]\[22\] _03768_
+ VGND VGND VPWR VPWR _03769_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_118_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09155_ net923 net4401 net575 VGND VGND VPWR VPWR _00909_ sky130_fd_sc_hd__mux2_1
XFILLER_166_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06367_ tag_array.tag0\[13\]\[16\] net1599 net1503 tag_array.tag0\[14\]\[16\] VGND
+ VGND VPWR VPWR _03706_ sky130_fd_sc_hd__a22o_1
XFILLER_135_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08106_ data_array.data1\[12\]\[60\] net1414 net1320 data_array.data1\[15\]\[60\]
+ _05286_ VGND VGND VPWR VPWR _05287_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_135_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09086_ net940 net3890 net416 VGND VGND VPWR VPWR _00840_ sky130_fd_sc_hd__mux2_1
X_06298_ tag_array.tag0\[12\]\[10\] net1405 net1311 tag_array.tag0\[15\]\[10\] _03642_
+ VGND VGND VPWR VPWR _03643_ sky130_fd_sc_hd__a221o_1
XFILLER_135_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08037_ data_array.data1\[1\]\[54\] net1544 net1448 data_array.data1\[2\]\[54\] VGND
+ VGND VPWR VPWR _05224_ sky130_fd_sc_hd__a22o_1
XFILLER_163_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold840 data_array.data1\[9\]\[36\] VGND VGND VPWR VPWR net2491 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold851 data_array.data1\[12\]\[31\] VGND VGND VPWR VPWR net2502 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold862 data_array.data0\[7\]\[10\] VGND VGND VPWR VPWR net2513 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold873 tag_array.tag1\[12\]\[5\] VGND VGND VPWR VPWR net2524 sky130_fd_sc_hd__dlygate4sd3_1
Xhold884 data_array.data0\[9\]\[60\] VGND VGND VPWR VPWR net2535 sky130_fd_sc_hd__dlygate4sd3_1
Xhold895 data_array.data1\[3\]\[30\] VGND VGND VPWR VPWR net2546 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_107_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09988_ net877 net2743 net372 VGND VGND VPWR VPWR _01737_ sky130_fd_sc_hd__mux2_1
XFILLER_130_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2230 data_array.data0\[15\]\[11\] VGND VGND VPWR VPWR net3881 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_114_1018 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2241 data_array.data1\[12\]\[43\] VGND VGND VPWR VPWR net3892 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2252 data_array.data0\[14\]\[30\] VGND VGND VPWR VPWR net3903 sky130_fd_sc_hd__dlygate4sd3_1
X_08939_ net1009 net2816 net426 VGND VGND VPWR VPWR _00695_ sky130_fd_sc_hd__mux2_1
Xhold2263 data_array.data0\[12\]\[63\] VGND VGND VPWR VPWR net3914 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2274 data_array.data1\[11\]\[36\] VGND VGND VPWR VPWR net3925 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_150_Right_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1540 data_array.data0\[8\]\[20\] VGND VGND VPWR VPWR net3191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2285 tag_array.tag1\[9\]\[14\] VGND VGND VPWR VPWR net3936 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1551 data_array.data1\[14\]\[46\] VGND VGND VPWR VPWR net3202 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2296 tag_array.tag1\[14\]\[19\] VGND VGND VPWR VPWR net3947 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1562 tag_array.tag1\[9\]\[13\] VGND VGND VPWR VPWR net3213 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11950_ clknet_leaf_92_clk _00758_ VGND VGND VPWR VPWR data_array.data0\[4\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1573 data_array.data0\[3\]\[5\] VGND VGND VPWR VPWR net3224 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_177_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1584 data_array.data0\[8\]\[58\] VGND VGND VPWR VPWR net3235 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_28_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10901_ net883 net4148 net514 VGND VGND VPWR VPWR _02646_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1595 lru_array.lru_mem\[4\] VGND VGND VPWR VPWR net3246 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_83_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_298 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11881_ clknet_leaf_58_clk _00689_ VGND VGND VPWR VPWR data_array.data0\[5\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13620_ clknet_leaf_22_clk _02249_ VGND VGND VPWR VPWR data_array.data0\[9\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
X_10832_ net2292 net900 net505 VGND VGND VPWR VPWR _02577_ sky130_fd_sc_hd__mux2_1
X_13551_ clknet_leaf_75_clk _02180_ VGND VGND VPWR VPWR data_array.data1\[0\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
X_10763_ net922 net4223 net498 VGND VGND VPWR VPWR _02508_ sky130_fd_sc_hd__mux2_1
X_12502_ clknet_leaf_216_clk _01196_ VGND VGND VPWR VPWR data_array.data1\[9\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13482_ clknet_leaf_145_clk _02112_ VGND VGND VPWR VPWR tag_array.tag0\[15\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_157_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10694_ net2912 net942 net485 VGND VGND VPWR VPWR _02439_ sky130_fd_sc_hd__mux2_1
XFILLER_139_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12433_ clknet_leaf_1_clk _01127_ VGND VGND VPWR VPWR data_array.data0\[14\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_139_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12364_ clknet_leaf_257_clk _00040_ VGND VGND VPWR VPWR data_array.rdata0\[46\] sky130_fd_sc_hd__dfxtp_1
X_14103_ clknet_leaf_63_clk _02732_ VGND VGND VPWR VPWR data_array.data0\[1\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_11315_ net1034 net3409 net801 VGND VGND VPWR VPWR _03058_ sky130_fd_sc_hd__mux2_1
XFILLER_5_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12295_ clknet_leaf_32_clk _01053_ VGND VGND VPWR VPWR tag_array.tag1\[12\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_14034_ clknet_leaf_116_clk _02663_ VGND VGND VPWR VPWR data_array.data1\[6\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11246_ net1045 net3206 net677 VGND VGND VPWR VPWR _02989_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11177_ net1066 net3292 net660 VGND VGND VPWR VPWR _02920_ sky130_fd_sc_hd__mux2_1
XFILLER_122_774 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10128_ net1032 net3279 net367 VGND VGND VPWR VPWR _01876_ sky130_fd_sc_hd__mux2_1
XFILLER_0_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10059_ net789 net2846 net599 VGND VGND VPWR VPWR _01808_ sky130_fd_sc_hd__mux2_1
XFILLER_76_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13818_ clknet_leaf_259_clk _02447_ VGND VGND VPWR VPWR data_array.data1\[2\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13749_ clknet_leaf_26_clk _02378_ VGND VGND VPWR VPWR data_array.data1\[1\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
X_07270_ data_array.data0\[12\]\[48\] net1391 net1297 data_array.data0\[15\]\[48\]
+ _04526_ VGND VGND VPWR VPWR _04527_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_14_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06221_ tag_array.tag0\[12\]\[3\] net1373 net1280 tag_array.tag0\[15\]\[3\] _03572_
+ VGND VGND VPWR VPWR _03573_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_152_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06152_ net27 net26 VGND VGND VPWR VPWR _03509_ sky130_fd_sc_hd__nand2b_2
XTAP_TAPCELL_ROW_152_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold103 data_array.data0\[8\]\[5\] VGND VGND VPWR VPWR net1754 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_866 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold114 tag_array.tag1\[8\]\[22\] VGND VGND VPWR VPWR net1765 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold125 data_array.data1\[1\]\[5\] VGND VGND VPWR VPWR net1776 sky130_fd_sc_hd__dlygate4sd3_1
X_06083_ net1159 net25 fsm.tag_out1\[24\] net1131 VGND VGND VPWR VPWR _03505_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_113_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold136 data_array.data1\[1\]\[13\] VGND VGND VPWR VPWR net1787 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_7_clk clknet_5_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_117_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold147 data_array.data1\[0\]\[7\] VGND VGND VPWR VPWR net1798 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold158 data_array.data0\[4\]\[9\] VGND VGND VPWR VPWR net1809 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09911_ net762 net4517 net604 VGND VGND VPWR VPWR _01661_ sky130_fd_sc_hd__mux2_1
Xhold169 data_array.data0\[0\]\[31\] VGND VGND VPWR VPWR net1820 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_99_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout605 net608 VGND VGND VPWR VPWR net605 sky130_fd_sc_hd__buf_4
Xfanout616 _05571_ VGND VGND VPWR VPWR net616 sky130_fd_sc_hd__buf_4
X_09842_ net1103 net2534 net380 VGND VGND VPWR VPWR _01592_ sky130_fd_sc_hd__mux2_1
XFILLER_86_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout627 net629 VGND VGND VPWR VPWR net627 sky130_fd_sc_hd__buf_4
Xfanout638 _05557_ VGND VGND VPWR VPWR net638 sky130_fd_sc_hd__clkbuf_8
XFILLER_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout649 net651 VGND VGND VPWR VPWR net649 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09773_ net1920 net695 net665 VGND VGND VPWR VPWR _01525_ sky130_fd_sc_hd__mux2_1
XFILLER_86_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06985_ data_array.data0\[5\]\[22\] net1533 net1437 data_array.data0\[6\]\[22\] VGND
+ VGND VPWR VPWR _04268_ sky130_fd_sc_hd__a22o_1
XFILLER_74_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Left_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08724_ net2279 net728 net475 VGND VGND VPWR VPWR _00483_ sky130_fd_sc_hd__mux2_1
XFILLER_37_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_05936_ data_array.rdata0\[35\] net846 net1142 VGND VGND VPWR VPWR _03418_ sky130_fd_sc_hd__o21a_1
XFILLER_160_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08655_ net2463 net703 net506 VGND VGND VPWR VPWR _00414_ sky130_fd_sc_hd__mux2_1
XFILLER_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05867_ data_array.rdata0\[12\] net1659 net1149 VGND VGND VPWR VPWR _03372_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_159_3416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_159_3427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07606_ data_array.data1\[9\]\[15\] net1584 net1488 data_array.data1\[10\]\[15\]
+ VGND VGND VPWR VPWR _04832_ sky130_fd_sc_hd__a22o_1
X_08586_ net780 net3845 net529 VGND VGND VPWR VPWR _00345_ sky130_fd_sc_hd__mux2_1
X_05798_ _03294_ _03303_ _03307_ _03314_ VGND VGND VPWR VPWR _03315_ sky130_fd_sc_hd__nor4_2
XTAP_TAPCELL_ROW_176_3741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07537_ net1192 _04763_ _04767_ net1618 VGND VGND VPWR VPWR _04770_ sky130_fd_sc_hd__a22o_1
XFILLER_23_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07468_ data_array.data1\[8\]\[2\] net1339 net1245 data_array.data1\[11\]\[2\] _04706_
+ VGND VGND VPWR VPWR _04707_ sky130_fd_sc_hd__a221o_1
XFILLER_139_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09207_ net752 net4436 net631 VGND VGND VPWR VPWR _00961_ sky130_fd_sc_hd__mux2_1
X_06419_ tag_array.tag0\[12\]\[21\] net1408 net1314 tag_array.tag0\[15\]\[21\] _03752_
+ VGND VGND VPWR VPWR _03753_ sky130_fd_sc_hd__a221o_1
XFILLER_120_1000 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07399_ data_array.data0\[5\]\[60\] net1603 net1507 data_array.data0\[6\]\[60\] VGND
+ VGND VPWR VPWR _04644_ sky130_fd_sc_hd__a22o_1
X_09138_ net991 net3732 net574 VGND VGND VPWR VPWR _00892_ sky130_fd_sc_hd__mux2_1
XFILLER_135_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09069_ net1009 net4198 net410 VGND VGND VPWR VPWR _00823_ sky130_fd_sc_hd__mux2_1
XFILLER_2_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11100_ net1763 net860 net335 VGND VGND VPWR VPWR _02843_ sky130_fd_sc_hd__mux2_1
XFILLER_162_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12080_ clknet_leaf_255_clk _00888_ VGND VGND VPWR VPWR data_array.data1\[14\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_150_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold670 tag_array.tag1\[6\]\[18\] VGND VGND VPWR VPWR net2321 sky130_fd_sc_hd__dlygate4sd3_1
Xhold681 data_array.data1\[7\]\[23\] VGND VGND VPWR VPWR net2332 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold692 tag_array.tag1\[15\]\[18\] VGND VGND VPWR VPWR net2343 sky130_fd_sc_hd__dlygate4sd3_1
X_11031_ net2500 net876 net338 VGND VGND VPWR VPWR _02775_ sky130_fd_sc_hd__mux2_1
XFILLER_104_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2060 data_array.data1\[5\]\[7\] VGND VGND VPWR VPWR net3711 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2071 data_array.data1\[5\]\[16\] VGND VGND VPWR VPWR net3722 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_134_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2082 tag_array.tag1\[9\]\[7\] VGND VGND VPWR VPWR net3733 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2093 data_array.data0\[3\]\[21\] VGND VGND VPWR VPWR net3744 sky130_fd_sc_hd__dlygate4sd3_1
X_12982_ clknet_leaf_182_clk _01676_ VGND VGND VPWR VPWR tag_array.tag0\[4\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_92_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1370 data_array.data0\[2\]\[48\] VGND VGND VPWR VPWR net3021 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1381 tag_array.tag1\[2\]\[9\] VGND VGND VPWR VPWR net3032 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11933_ clknet_leaf_112_clk _00741_ VGND VGND VPWR VPWR data_array.data0\[4\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1392 data_array.data1\[13\]\[26\] VGND VGND VPWR VPWR net3043 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11864_ clknet_leaf_247_clk _00672_ VGND VGND VPWR VPWR data_array.data0\[5\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13603_ clknet_leaf_31_clk _02232_ VGND VGND VPWR VPWR data_array.data0\[9\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_10815_ net4280 net968 net504 VGND VGND VPWR VPWR _02560_ sky130_fd_sc_hd__mux2_1
X_11795_ clknet_leaf_192_clk _00603_ VGND VGND VPWR VPWR data_array.data0\[8\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13534_ clknet_leaf_44_clk _02163_ VGND VGND VPWR VPWR data_array.data1\[0\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_10746_ net990 net2546 net497 VGND VGND VPWR VPWR _02491_ sky130_fd_sc_hd__mux2_1
XFILLER_14_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13465_ clknet_leaf_162_clk _02095_ VGND VGND VPWR VPWR tag_array.tag0\[1\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_10677_ net2839 net1008 net478 VGND VGND VPWR VPWR _02422_ sky130_fd_sc_hd__mux2_1
X_12416_ clknet_leaf_11_clk _01110_ VGND VGND VPWR VPWR data_array.data0\[14\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_173_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13396_ clknet_leaf_213_clk _02026_ VGND VGND VPWR VPWR data_array.data1\[8\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_58_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput208 net208 VGND VGND VPWR VPWR cpu_rdata[49] sky130_fd_sc_hd__buf_6
XFILLER_57_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12347_ clknet_leaf_52_clk _00021_ VGND VGND VPWR VPWR data_array.rdata0\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_153_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput219 net219 VGND VGND VPWR VPWR cpu_rdata[59] sky130_fd_sc_hd__clkbuf_4
XFILLER_126_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_387 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12278_ clknet_leaf_105_clk _01036_ VGND VGND VPWR VPWR tag_array.tag1\[13\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_49_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14017_ clknet_leaf_249_clk _02646_ VGND VGND VPWR VPWR data_array.data1\[5\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11229_ net859 net3559 net652 VGND VGND VPWR VPWR _02972_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_711 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06770_ data_array.data0\[13\]\[3\] net1567 net1471 data_array.data0\[14\]\[3\] VGND
+ VGND VPWR VPWR _04072_ sky130_fd_sc_hd__a22o_1
XFILLER_49_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05721_ net22 fsm.tag_out1\[22\] VGND VGND VPWR VPWR _03238_ sky130_fd_sc_hd__xor2_1
XFILLER_36_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08440_ net1124 _05529_ VGND VGND VPWR VPWR _05530_ sky130_fd_sc_hd__and2_1
X_05652_ net3 fsm.tag_out0\[4\] VGND VGND VPWR VPWR _03169_ sky130_fd_sc_hd__and2b_1
XFILLER_56_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08371_ net1123 _05483_ VGND VGND VPWR VPWR _05484_ sky130_fd_sc_hd__and2_1
XFILLER_56_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07322_ data_array.data0\[1\]\[53\] net1524 net1428 data_array.data0\[2\]\[53\] VGND
+ VGND VPWR VPWR _04574_ sky130_fd_sc_hd__a22o_1
XFILLER_143_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_945 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07253_ _04510_ _04511_ VGND VGND VPWR VPWR _00040_ sky130_fd_sc_hd__or2_1
XFILLER_104_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06204_ tag_array.tag0\[1\]\[1\] net1592 net1496 tag_array.tag0\[2\]\[1\] VGND VGND
+ VPWR VPWR _03558_ sky130_fd_sc_hd__a22o_1
X_07184_ data_array.data0\[0\]\[40\] net1412 net1318 data_array.data0\[3\]\[40\] _04448_
+ VGND VGND VPWR VPWR _04449_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_132_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06135_ data_array.rdata0\[50\] net1135 net1116 data_array.rdata1\[50\] VGND VGND
+ VPWR VPWR net308 sky130_fd_sc_hd__a22o_1
XFILLER_2_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06066_ fsm.tag_out0\[15\] net1122 _03496_ VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__a21o_1
Xfanout402 net403 VGND VGND VPWR VPWR net402 sky130_fd_sc_hd__buf_4
XFILLER_160_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout413 net417 VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__buf_4
XFILLER_59_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout424 net425 VGND VGND VPWR VPWR net424 sky130_fd_sc_hd__buf_4
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Left_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout435 net441 VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__clkbuf_4
Xfanout446 net448 VGND VGND VPWR VPWR net446 sky130_fd_sc_hd__clkbuf_8
XFILLER_141_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout457 net458 VGND VGND VPWR VPWR net457 sky130_fd_sc_hd__buf_4
X_09825_ net909 net3259 net387 VGND VGND VPWR VPWR _01576_ sky130_fd_sc_hd__mux2_1
Xfanout468 net477 VGND VGND VPWR VPWR net468 sky130_fd_sc_hd__buf_4
XFILLER_171_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout479 net480 VGND VGND VPWR VPWR net479 sky130_fd_sc_hd__clkbuf_8
X_09756_ net2565 net764 net671 VGND VGND VPWR VPWR _01508_ sky130_fd_sc_hd__mux2_1
X_06968_ data_array.data0\[9\]\[21\] net1555 net1459 data_array.data0\[10\]\[21\]
+ VGND VGND VPWR VPWR _04252_ sky130_fd_sc_hd__a22o_1
XFILLER_73_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08707_ net2290 net694 net482 VGND VGND VPWR VPWR _00466_ sky130_fd_sc_hd__mux2_1
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05919_ data_array.rdata1\[29\] net833 net842 VGND VGND VPWR VPWR _03407_ sky130_fd_sc_hd__a21o_1
X_09687_ net738 net3798 net606 VGND VGND VPWR VPWR _01439_ sky130_fd_sc_hd__mux2_1
X_06899_ net1628 _04183_ _04187_ net1202 VGND VGND VPWR VPWR _04190_ sky130_fd_sc_hd__a22o_1
XFILLER_55_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08638_ net2344 net773 net510 VGND VGND VPWR VPWR _00397_ sky130_fd_sc_hd__mux2_1
XFILLER_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_10 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08569_ net811 _05577_ net1698 VGND VGND VPWR VPWR _00335_ sky130_fd_sc_hd__a21o_1
XFILLER_70_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_30_Left_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10600_ net2117 net1062 net472 VGND VGND VPWR VPWR _02345_ sky130_fd_sc_hd__mux2_1
XFILLER_11_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11580_ clknet_leaf_100_clk _00388_ VGND VGND VPWR VPWR tag_array.tag1\[5\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_10531_ net1083 net2693 net462 VGND VGND VPWR VPWR _02276_ sky130_fd_sc_hd__mux2_1
XFILLER_7_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire836 _03315_ VGND VGND VPWR VPWR net836 sky130_fd_sc_hd__buf_2
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13250_ clknet_leaf_176_clk _01880_ VGND VGND VPWR VPWR data_array.data0\[11\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_10462_ net1096 net3261 net348 VGND VGND VPWR VPWR _02207_ sky130_fd_sc_hd__mux2_1
XFILLER_10_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12201_ clknet_leaf_148_clk _00154_ VGND VGND VPWR VPWR fsm.tag_out0\[8\] sky130_fd_sc_hd__dfxtp_1
X_13181_ clknet_leaf_15_clk _00073_ VGND VGND VPWR VPWR data_array.rdata1\[18\] sky130_fd_sc_hd__dfxtp_1
X_10393_ net1798 net1083 net668 VGND VGND VPWR VPWR _02139_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_92_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12132_ clknet_leaf_171_clk _00940_ VGND VGND VPWR VPWR tag_array.tag0\[12\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12063_ clknet_leaf_57_clk _00871_ VGND VGND VPWR VPWR data_array.data1\[14\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11014_ net1965 net946 net336 VGND VGND VPWR VPWR _02758_ sky130_fd_sc_hd__mux2_1
XFILLER_49_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout980 _05484_ VGND VGND VPWR VPWR net980 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_240_clk clknet_5_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_240_clk
+ sky130_fd_sc_hd__clkbuf_8
Xfanout991 _05480_ VGND VGND VPWR VPWR net991 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_5_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12965_ clknet_leaf_143_clk _01659_ VGND VGND VPWR VPWR tag_array.tag0\[4\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_11916_ clknet_leaf_221_clk _00724_ VGND VGND VPWR VPWR data_array.data0\[5\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_16_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12896_ clknet_leaf_230_clk _01590_ VGND VGND VPWR VPWR data_array.data0\[13\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_11847_ clknet_leaf_53_clk _00655_ VGND VGND VPWR VPWR data_array.data0\[7\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_159_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11778_ clknet_leaf_84_clk _00586_ VGND VGND VPWR VPWR data_array.data0\[8\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_159_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13517_ clknet_leaf_42_clk _02146_ VGND VGND VPWR VPWR data_array.data1\[0\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_158_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10729_ net1056 net3192 net493 VGND VGND VPWR VPWR _02474_ sky130_fd_sc_hd__mux2_1
X_14497_ clknet_leaf_171_clk _00129_ VGND VGND VPWR VPWR dirty_way0 sky130_fd_sc_hd__dfxtp_1
Xclkload12 clknet_5_27__leaf_clk VGND VGND VPWR VPWR clkload12/Y sky130_fd_sc_hd__inv_6
XFILLER_16_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13448_ clknet_leaf_191_clk _02078_ VGND VGND VPWR VPWR tag_array.tag0\[1\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload23 clknet_leaf_262_clk VGND VGND VPWR VPWR clkload23/Y sky130_fd_sc_hd__inv_6
Xclkload34 clknet_leaf_15_clk VGND VGND VPWR VPWR clkload34/Y sky130_fd_sc_hd__bufinv_16
Xclkload45 clknet_leaf_245_clk VGND VGND VPWR VPWR clkload45/Y sky130_fd_sc_hd__clkinv_4
Xclkload56 clknet_leaf_254_clk VGND VGND VPWR VPWR clkload56/X sky130_fd_sc_hd__clkbuf_8
XFILLER_103_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13379_ clknet_leaf_190_clk _02009_ VGND VGND VPWR VPWR tag_array.tag0\[2\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload67 clknet_leaf_31_clk VGND VGND VPWR VPWR clkload67/Y sky130_fd_sc_hd__bufinv_16
Xclkload78 clknet_leaf_50_clk VGND VGND VPWR VPWR clkload78/Y sky130_fd_sc_hd__inv_6
XFILLER_127_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload89 clknet_leaf_61_clk VGND VGND VPWR VPWR clkload89/X sky130_fd_sc_hd__clkbuf_4
XFILLER_69_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07940_ data_array.data1\[9\]\[45\] net1540 net1444 data_array.data1\[10\]\[45\]
+ VGND VGND VPWR VPWR _05136_ sky130_fd_sc_hd__a22o_1
Xhold2807 tag_array.dirty1\[7\] VGND VGND VPWR VPWR net4458 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_142_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2818 tag_array.tag0\[12\]\[17\] VGND VGND VPWR VPWR net4469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2829 data_array.data0\[3\]\[56\] VGND VGND VPWR VPWR net4480 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_147_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07871_ data_array.data1\[8\]\[39\] net1347 net1253 data_array.data1\[11\]\[39\]
+ _05072_ VGND VGND VPWR VPWR _05073_ sky130_fd_sc_hd__a221o_1
XFILLER_110_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_147_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09610_ net909 net4428 net395 VGND VGND VPWR VPWR _01362_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_231_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_231_clk
+ sky130_fd_sc_hd__clkbuf_8
X_06822_ net1631 _04113_ _04117_ net1205 VGND VGND VPWR VPWR _04120_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_108_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09541_ net763 net3703 net620 VGND VGND VPWR VPWR _01294_ sky130_fd_sc_hd__mux2_1
X_06753_ data_array.data0\[8\]\[1\] net1333 net1239 data_array.data0\[11\]\[1\] _04056_
+ VGND VGND VPWR VPWR _04057_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_125_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05704_ net30 fsm.tag_out0\[0\] VGND VGND VPWR VPWR _03221_ sky130_fd_sc_hd__or2_1
X_09472_ net741 net3872 net659 VGND VGND VPWR VPWR _01225_ sky130_fd_sc_hd__mux2_1
XFILLER_52_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06684_ tag_array.tag1\[1\]\[20\] net1541 net1445 tag_array.tag1\[2\]\[20\] VGND
+ VGND VPWR VPWR _03994_ sky130_fd_sc_hd__a22o_1
XFILLER_34_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08423_ net1750 net912 net691 VGND VGND VPWR VPWR _00270_ sky130_fd_sc_hd__mux2_1
XFILLER_169_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05635_ _03134_ net4626 _03150_ net4625 VGND VGND VPWR VPWR _00187_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_121_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08354_ net2512 net1007 net689 VGND VGND VPWR VPWR _00247_ sky130_fd_sc_hd__mux2_1
XFILLER_177_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07305_ data_array.data0\[0\]\[51\] net1332 net1238 data_array.data0\[3\]\[51\] _04558_
+ VGND VGND VPWR VPWR _04559_ sky130_fd_sc_hd__a221o_1
XFILLER_20_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08285_ net2266 net1096 net692 VGND VGND VPWR VPWR _00224_ sky130_fd_sc_hd__mux2_1
Xclkload6 clknet_5_12__leaf_clk VGND VGND VPWR VPWR clkload6/Y sky130_fd_sc_hd__inv_6
XFILLER_164_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07236_ data_array.data0\[9\]\[45\] net1533 net1437 data_array.data0\[10\]\[45\]
+ VGND VGND VPWR VPWR _04496_ sky130_fd_sc_hd__a22o_1
XFILLER_164_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07167_ data_array.data0\[8\]\[39\] net1349 net1255 data_array.data0\[11\]\[39\]
+ _04432_ VGND VGND VPWR VPWR _04433_ sky130_fd_sc_hd__a221o_1
XFILLER_133_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06118_ data_array.rdata0\[33\] net1139 net1115 data_array.rdata1\[33\] VGND VGND
+ VPWR VPWR net289 sky130_fd_sc_hd__a22o_1
X_07098_ net1214 _04365_ _04369_ net1165 VGND VGND VPWR VPWR _04371_ sky130_fd_sc_hd__a22o_1
XFILLER_106_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06049_ net1164 net6 fsm.tag_out1\[7\] net1132 VGND VGND VPWR VPWR _03488_ sky130_fd_sc_hd__a22o_1
Xfanout1208 net1211 VGND VGND VPWR VPWR net1208 sky130_fd_sc_hd__buf_4
XFILLER_121_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1219 net1220 VGND VGND VPWR VPWR net1219 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_184_3895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_222_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_222_clk
+ sky130_fd_sc_hd__clkbuf_8
X_09808_ net977 net3297 net391 VGND VGND VPWR VPWR _01559_ sky130_fd_sc_hd__mux2_1
XFILLER_28_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_105_Left_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_447 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09739_ net731 net4418 net680 VGND VGND VPWR VPWR _01491_ sky130_fd_sc_hd__mux2_1
XFILLER_28_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12750_ clknet_leaf_153_clk _01444_ VGND VGND VPWR VPWR tag_array.tag0\[5\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_131_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11701_ clknet_leaf_141_clk _00509_ VGND VGND VPWR VPWR tag_array.tag1\[15\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12681_ clknet_leaf_225_clk _01375_ VGND VGND VPWR VPWR data_array.data0\[15\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_43_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14420_ clknet_leaf_69_clk _03043_ VGND VGND VPWR VPWR data_array.data1\[7\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_11632_ clknet_leaf_129_clk _00440_ VGND VGND VPWR VPWR tag_array.tag1\[3\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_46_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_917 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14351_ clknet_leaf_265_clk _02974_ VGND VGND VPWR VPWR data_array.data1\[10\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_126_1072 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11563_ clknet_leaf_193_clk _00371_ VGND VGND VPWR VPWR tag_array.tag1\[5\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13302_ clknet_leaf_45_clk _01932_ VGND VGND VPWR VPWR data_array.data0\[10\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_42_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10514_ net889 net4506 net345 VGND VGND VPWR VPWR _02259_ sky130_fd_sc_hd__mux2_1
X_14282_ clknet_leaf_251_clk _02911_ VGND VGND VPWR VPWR data_array.data1\[11\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_11494_ clknet_leaf_153_clk _00303_ VGND VGND VPWR VPWR tag_array.valid0\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_21_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13233_ clknet_leaf_0_clk _01863_ VGND VGND VPWR VPWR data_array.data0\[11\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_170_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10445_ net1969 net874 net667 VGND VGND VPWR VPWR _02191_ sky130_fd_sc_hd__mux2_1
XFILLER_40_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13164_ clknet_leaf_266_clk _00075_ VGND VGND VPWR VPWR data_array.rdata1\[1\] sky130_fd_sc_hd__dfxtp_1
X_10376_ net696 net3366 net540 VGND VGND VPWR VPWR _02123_ sky130_fd_sc_hd__mux2_1
XFILLER_123_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12115_ clknet_leaf_210_clk _00923_ VGND VGND VPWR VPWR data_array.data1\[14\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_123_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13095_ clknet_leaf_6_clk _01789_ VGND VGND VPWR VPWR data_array.data1\[13\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_111_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12046_ clknet_leaf_12_clk _00854_ VGND VGND VPWR VPWR data_array.data0\[6\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_49_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_213_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_213_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_77_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13997_ clknet_leaf_215_clk _02626_ VGND VGND VPWR VPWR data_array.data1\[5\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_142_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12948_ clknet_leaf_224_clk _01642_ VGND VGND VPWR VPWR data_array.data0\[13\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12879_ clknet_leaf_38_clk _01573_ VGND VGND VPWR VPWR data_array.data0\[12\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_83_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_747 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08070_ data_array.data1\[1\]\[57\] net1528 net1432 data_array.data1\[2\]\[57\] VGND
+ VGND VPWR VPWR _05254_ sky130_fd_sc_hd__a22o_1
XFILLER_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload101 clknet_leaf_36_clk VGND VGND VPWR VPWR clkload101/X sky130_fd_sc_hd__clkbuf_8
Xclkload112 clknet_leaf_95_clk VGND VGND VPWR VPWR clkload112/Y sky130_fd_sc_hd__inv_8
Xclkload123 clknet_leaf_78_clk VGND VGND VPWR VPWR clkload123/Y sky130_fd_sc_hd__inv_6
XFILLER_128_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload134 clknet_leaf_216_clk VGND VGND VPWR VPWR clkload134/Y sky130_fd_sc_hd__inv_6
X_07021_ net1213 _04295_ _04299_ net1165 VGND VGND VPWR VPWR _04301_ sky130_fd_sc_hd__a22o_1
Xclkload145 clknet_leaf_210_clk VGND VGND VPWR VPWR clkload145/Y sky130_fd_sc_hd__clkinv_4
Xclkload156 clknet_leaf_169_clk VGND VGND VPWR VPWR clkload156/Y sky130_fd_sc_hd__bufinv_16
Xclkload167 clknet_leaf_205_clk VGND VGND VPWR VPWR clkload167/Y sky130_fd_sc_hd__inv_6
Xclkload178 clknet_leaf_178_clk VGND VGND VPWR VPWR clkload178/Y sky130_fd_sc_hd__clkinv_4
Xclkload189 clknet_leaf_190_clk VGND VGND VPWR VPWR clkload189/Y sky130_fd_sc_hd__inv_8
XFILLER_143_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08972_ net876 net2715 net429 VGND VGND VPWR VPWR _00728_ sky130_fd_sc_hd__mux2_1
Xhold2604 data_array.data0\[10\]\[48\] VGND VGND VPWR VPWR net4255 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2615 tag_array.tag1\[10\]\[19\] VGND VGND VPWR VPWR net4266 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2626 data_array.data0\[9\]\[56\] VGND VGND VPWR VPWR net4277 sky130_fd_sc_hd__dlygate4sd3_1
X_07923_ net1224 _05115_ _05119_ net1176 VGND VGND VPWR VPWR _05121_ sky130_fd_sc_hd__a22o_1
Xhold2637 data_array.data1\[6\]\[10\] VGND VGND VPWR VPWR net4288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2648 data_array.data1\[11\]\[25\] VGND VGND VPWR VPWR net4299 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1903 data_array.data0\[3\]\[0\] VGND VGND VPWR VPWR net3554 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1914 data_array.data1\[11\]\[20\] VGND VGND VPWR VPWR net3565 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_204_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_204_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold2659 data_array.data0\[8\]\[23\] VGND VGND VPWR VPWR net4310 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_127_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1925 tag_array.tag0\[8\]\[23\] VGND VGND VPWR VPWR net3576 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_162_3467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07854_ data_array.data1\[5\]\[37\] net1544 net1448 data_array.data1\[6\]\[37\] VGND
+ VGND VPWR VPWR _05058_ sky130_fd_sc_hd__a22o_1
Xhold1936 tag_array.tag0\[1\]\[11\] VGND VGND VPWR VPWR net3587 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1947 data_array.data1\[8\]\[0\] VGND VGND VPWR VPWR net3598 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_162_3478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1958 data_array.data1\[6\]\[0\] VGND VGND VPWR VPWR net3609 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1969 data_array.data0\[3\]\[1\] VGND VGND VPWR VPWR net3620 sky130_fd_sc_hd__dlygate4sd3_1
X_06805_ data_array.data0\[1\]\[6\] net1519 net1423 data_array.data0\[2\]\[6\] VGND
+ VGND VPWR VPWR _04104_ sky130_fd_sc_hd__a22o_1
XFILLER_44_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07785_ data_array.data1\[4\]\[31\] net1381 net1287 data_array.data1\[7\]\[31\] _04994_
+ VGND VGND VPWR VPWR _04995_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_123_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09524_ net733 net2408 net622 VGND VGND VPWR VPWR _01277_ sky130_fd_sc_hd__mux2_1
X_06736_ _04040_ _04041_ VGND VGND VPWR VPWR _00172_ sky130_fd_sc_hd__or2_1
X_09455_ net819 net3481 _05596_ VGND VGND VPWR VPWR _01208_ sky130_fd_sc_hd__mux2_1
XFILLER_169_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06667_ tag_array.tag1\[4\]\[18\] net1372 net1278 tag_array.tag1\[7\]\[18\] _03978_
+ VGND VGND VPWR VPWR _03979_ sky130_fd_sc_hd__a221o_1
XFILLER_101_34 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08406_ net137 net72 net1642 VGND VGND VPWR VPWR _05507_ sky130_fd_sc_hd__mux2_1
XFILLER_52_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05618_ net14 VGND VGND VPWR VPWR _03140_ sky130_fd_sc_hd__inv_2
X_09386_ net857 net3934 net404 VGND VGND VPWR VPWR _01139_ sky130_fd_sc_hd__mux2_1
X_06598_ tag_array.tag1\[9\]\[12\] net1592 net1496 tag_array.tag1\[10\]\[12\] VGND
+ VGND VPWR VPWR _03916_ sky130_fd_sc_hd__a22o_1
XFILLER_177_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08337_ net112 net47 net1643 VGND VGND VPWR VPWR _05461_ sky130_fd_sc_hd__mux2_1
XFILLER_131_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08268_ net694 net3500 net799 VGND VGND VPWR VPWR _00220_ sky130_fd_sc_hd__mux2_1
XFILLER_137_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_705 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07219_ net1224 _04475_ _04479_ net1176 VGND VGND VPWR VPWR _04481_ sky130_fd_sc_hd__a22o_1
X_08199_ net787 net4211 net805 VGND VGND VPWR VPWR _00197_ sky130_fd_sc_hd__mux2_1
X_10230_ net884 net3735 net354 VGND VGND VPWR VPWR _01977_ sky130_fd_sc_hd__mux2_1
XFILLER_105_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_750 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_964 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10161_ net902 net2723 net364 VGND VGND VPWR VPWR _01909_ sky130_fd_sc_hd__mux2_1
XFILLER_0_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1005 _05472_ VGND VGND VPWR VPWR net1005 sky130_fd_sc_hd__clkbuf_2
Xfanout1016 _05466_ VGND VGND VPWR VPWR net1016 sky130_fd_sc_hd__clkbuf_2
Xfanout1027 _05462_ VGND VGND VPWR VPWR net1027 sky130_fd_sc_hd__clkbuf_2
XFILLER_121_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10092_ net2740 net757 net642 VGND VGND VPWR VPWR _01841_ sky130_fd_sc_hd__mux2_1
Xfanout1038 _05456_ VGND VGND VPWR VPWR net1038 sky130_fd_sc_hd__clkbuf_2
XFILLER_121_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1049 net1051 VGND VGND VPWR VPWR net1049 sky130_fd_sc_hd__clkbuf_2
XFILLER_102_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13920_ clknet_leaf_93_clk _02549_ VGND VGND VPWR VPWR data_array.data1\[4\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13851_ clknet_leaf_66_clk _02480_ VGND VGND VPWR VPWR data_array.data1\[3\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_87_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12802_ clknet_leaf_231_clk _01496_ VGND VGND VPWR VPWR tag_array.tag1\[10\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_48_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13782_ clknet_leaf_47_clk _02411_ VGND VGND VPWR VPWR data_array.data1\[2\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_10994_ net1935 net1027 net339 VGND VGND VPWR VPWR _02738_ sky130_fd_sc_hd__mux2_1
XFILLER_16_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12733_ clknet_leaf_164_clk _01427_ VGND VGND VPWR VPWR tag_array.tag0\[5\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ clknet_leaf_23_clk _01358_ VGND VGND VPWR VPWR data_array.data0\[15\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_26_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_861 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14403_ clknet_leaf_5_clk _03026_ VGND VGND VPWR VPWR data_array.data1\[10\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
X_11615_ clknet_leaf_189_clk _00423_ VGND VGND VPWR VPWR tag_array.tag1\[3\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_61_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12595_ clknet_leaf_168_clk _01289_ VGND VGND VPWR VPWR tag_array.tag0\[0\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14334_ clknet_leaf_216_clk _02963_ VGND VGND VPWR VPWR data_array.data1\[11\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11546_ clknet_leaf_166_clk _00354_ VGND VGND VPWR VPWR tag_array.tag1\[6\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_171_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14265_ clknet_leaf_56_clk _02894_ VGND VGND VPWR VPWR data_array.data1\[12\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_167_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11477_ clknet_leaf_172_clk _00287_ VGND VGND VPWR VPWR tag_array.valid1\[11\] sky130_fd_sc_hd__dfxtp_1
X_13216_ clknet_leaf_2_clk _00112_ VGND VGND VPWR VPWR data_array.rdata1\[53\] sky130_fd_sc_hd__dfxtp_1
X_10428_ net2319 net942 net669 VGND VGND VPWR VPWR _02174_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_164_Right_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14196_ clknet_leaf_87_clk _02825_ VGND VGND VPWR VPWR data_array.data0\[2\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
X_13147_ clknet_leaf_142_clk _01841_ VGND VGND VPWR VPWR tag_array.tag1\[8\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_10359_ net762 net2727 net540 VGND VGND VPWR VPWR _02106_ sky130_fd_sc_hd__mux2_1
XFILLER_183_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13078_ clknet_leaf_39_clk _01772_ VGND VGND VPWR VPWR data_array.data1\[13\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_144_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1550 net1551 VGND VGND VPWR VPWR net1550 sky130_fd_sc_hd__clkbuf_4
X_12029_ clknet_leaf_241_clk _00837_ VGND VGND VPWR VPWR data_array.data0\[6\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_144_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1561 net1563 VGND VGND VPWR VPWR net1561 sky130_fd_sc_hd__clkbuf_4
XFILLER_93_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1572 net1573 VGND VGND VPWR VPWR net1572 sky130_fd_sc_hd__clkbuf_4
Xfanout1583 net1584 VGND VGND VPWR VPWR net1583 sky130_fd_sc_hd__clkbuf_4
XFILLER_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1594 net1613 VGND VGND VPWR VPWR net1594 sky130_fd_sc_hd__buf_2
XFILLER_54_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07570_ net1629 _04793_ _04797_ net1203 VGND VGND VPWR VPWR _04800_ sky130_fd_sc_hd__a22o_1
XFILLER_80_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06521_ tag_array.tag1\[13\]\[5\] net1608 net1512 tag_array.tag1\[14\]\[5\] VGND
+ VGND VPWR VPWR _03846_ sky130_fd_sc_hd__a22o_1
XFILLER_33_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09240_ net720 net3623 net645 VGND VGND VPWR VPWR _00994_ sky130_fd_sc_hd__mux2_1
X_06452_ tag_array.tag0\[8\]\[24\] net1374 net1281 tag_array.tag0\[11\]\[24\] _03782_
+ VGND VGND VPWR VPWR _03783_ sky130_fd_sc_hd__a221o_1
XFILLER_61_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09171_ net859 net2849 net570 VGND VGND VPWR VPWR _00925_ sky130_fd_sc_hd__mux2_1
X_06383_ net1183 _03715_ _03719_ net1231 VGND VGND VPWR VPWR _03721_ sky130_fd_sc_hd__a22o_1
X_08122_ _05300_ _05301_ VGND VGND VPWR VPWR _00121_ sky130_fd_sc_hd__or2_1
XFILLER_179_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08053_ data_array.data1\[4\]\[55\] net1343 net1249 data_array.data1\[7\]\[55\] _05238_
+ VGND VGND VPWR VPWR _05239_ sky130_fd_sc_hd__a221o_1
XFILLER_179_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07004_ data_array.data0\[4\]\[24\] net1386 net1292 data_array.data0\[7\]\[24\] _04284_
+ VGND VGND VPWR VPWR _04285_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_116_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_131_Right_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_164_3507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_102 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2401 data_array.data1\[10\]\[39\] VGND VGND VPWR VPWR net4052 sky130_fd_sc_hd__dlygate4sd3_1
X_08955_ net946 net4095 net426 VGND VGND VPWR VPWR _00711_ sky130_fd_sc_hd__mux2_1
Xinput108 mem_rdata[18] VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_1
Xhold2412 data_array.data0\[15\]\[28\] VGND VGND VPWR VPWR net4063 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_181_3832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2423 data_array.data0\[5\]\[16\] VGND VGND VPWR VPWR net4074 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput119 mem_rdata[28] VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_181_3843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2434 data_array.data0\[7\]\[59\] VGND VGND VPWR VPWR net4085 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2445 data_array.data1\[6\]\[39\] VGND VGND VPWR VPWR net4096 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1700 data_array.data0\[10\]\[42\] VGND VGND VPWR VPWR net3351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1711 data_array.data1\[13\]\[58\] VGND VGND VPWR VPWR net3362 sky130_fd_sc_hd__dlygate4sd3_1
X_07906_ data_array.data1\[4\]\[42\] net1399 net1305 data_array.data1\[7\]\[42\] _05104_
+ VGND VGND VPWR VPWR _05105_ sky130_fd_sc_hd__a221o_1
Xhold2456 data_array.data0\[13\]\[54\] VGND VGND VPWR VPWR net4107 sky130_fd_sc_hd__dlygate4sd3_1
X_08886_ net961 net2407 net436 VGND VGND VPWR VPWR _00643_ sky130_fd_sc_hd__mux2_1
Xhold1722 lru_array.lru_mem\[5\] VGND VGND VPWR VPWR net3373 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2467 tag_array.tag0\[0\]\[2\] VGND VGND VPWR VPWR net4118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1733 data_array.data1\[11\]\[40\] VGND VGND VPWR VPWR net3384 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2478 data_array.data0\[14\]\[57\] VGND VGND VPWR VPWR net4129 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2489 tag_array.tag1\[13\]\[12\] VGND VGND VPWR VPWR net4140 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1744 tag_array.tag0\[10\]\[8\] VGND VGND VPWR VPWR net3395 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1755 data_array.data1\[10\]\[55\] VGND VGND VPWR VPWR net3406 sky130_fd_sc_hd__dlygate4sd3_1
X_07837_ data_array.data1\[9\]\[36\] net1606 net1510 data_array.data1\[10\]\[36\]
+ VGND VGND VPWR VPWR _05042_ sky130_fd_sc_hd__a22o_1
Xhold1766 data_array.data0\[12\]\[13\] VGND VGND VPWR VPWR net3417 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1777 data_array.data1\[9\]\[54\] VGND VGND VPWR VPWR net3428 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_99_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1788 tag_array.tag0\[4\]\[19\] VGND VGND VPWR VPWR net3439 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1799 tag_array.tag0\[9\]\[18\] VGND VGND VPWR VPWR net3450 sky130_fd_sc_hd__dlygate4sd3_1
X_07768_ net1202 _04973_ _04977_ net1628 VGND VGND VPWR VPWR _04980_ sky130_fd_sc_hd__a22o_1
XFILLER_147_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09507_ net698 net4104 net625 VGND VGND VPWR VPWR _01260_ sky130_fd_sc_hd__mux2_1
X_06719_ tag_array.tag1\[13\]\[23\] net1610 net1514 tag_array.tag1\[14\]\[23\] VGND
+ VGND VPWR VPWR _04026_ sky130_fd_sc_hd__a22o_1
XFILLER_53_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_179_3794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07699_ data_array.data1\[8\]\[23\] net1361 net1267 data_array.data1\[11\]\[23\]
+ _04916_ VGND VGND VPWR VPWR _04917_ sky130_fd_sc_hd__a221o_1
X_09438_ net914 net3531 net585 VGND VGND VPWR VPWR _01191_ sky130_fd_sc_hd__mux2_1
XFILLER_169_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09369_ net926 net2441 net402 VGND VGND VPWR VPWR _01122_ sky130_fd_sc_hd__mux2_1
XFILLER_8_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11400_ clknet_leaf_232_clk _00210_ VGND VGND VPWR VPWR tag_array.tag1\[7\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_12380_ clknet_leaf_119_clk _00058_ VGND VGND VPWR VPWR data_array.rdata0\[62\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_70 _00039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_81 net520 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11331_ net968 net3383 net797 VGND VGND VPWR VPWR _03074_ sky130_fd_sc_hd__mux2_1
XANTENNA_92 net1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14050_ clknet_leaf_256_clk _02679_ VGND VGND VPWR VPWR data_array.data1\[6\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_11262_ net981 net4258 net673 VGND VGND VPWR VPWR _03005_ sky130_fd_sc_hd__mux2_1
XFILLER_181_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13001_ clknet_leaf_222_clk _01695_ VGND VGND VPWR VPWR data_array.data0\[3\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_10213_ net954 net3029 net355 VGND VGND VPWR VPWR _01960_ sky130_fd_sc_hd__mux2_1
X_11193_ net1001 net3764 net649 VGND VGND VPWR VPWR _02936_ sky130_fd_sc_hd__mux2_1
XFILLER_0_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10144_ net970 net2552 net363 VGND VGND VPWR VPWR _01892_ sky130_fd_sc_hd__mux2_1
XFILLER_67_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10075_ net722 net3562 net600 VGND VGND VPWR VPWR _01824_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_85_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1024 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13903_ clknet_leaf_82_clk _02532_ VGND VGND VPWR VPWR data_array.data1\[4\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_85_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13834_ clknet_leaf_251_clk _02463_ VGND VGND VPWR VPWR data_array.data1\[3\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13765_ clknet_leaf_211_clk _02394_ VGND VGND VPWR VPWR data_array.data1\[1\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_100_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10977_ net2838 net1092 net341 VGND VGND VPWR VPWR _02721_ sky130_fd_sc_hd__mux2_1
X_12716_ clknet_leaf_160_clk _01410_ VGND VGND VPWR VPWR tag_array.tag0\[7\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_13696_ clknet_leaf_21_clk _02325_ VGND VGND VPWR VPWR data_array.data1\[15\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_175_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12647_ clknet_leaf_55_clk _01341_ VGND VGND VPWR VPWR data_array.data0\[15\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_157_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12578_ clknet_leaf_107_clk _01272_ VGND VGND VPWR VPWR tag_array.tag0\[10\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14317_ clknet_leaf_213_clk _02946_ VGND VGND VPWR VPWR data_array.data1\[11\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
X_11529_ clknet_leaf_175_clk _00337_ VGND VGND VPWR VPWR tag_array.valid1\[3\] sky130_fd_sc_hd__dfxtp_1
Xhold307 data_array.data0\[6\]\[36\] VGND VGND VPWR VPWR net1958 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold318 data_array.data1\[0\]\[59\] VGND VGND VPWR VPWR net1969 sky130_fd_sc_hd__dlygate4sd3_1
Xhold329 data_array.data1\[8\]\[7\] VGND VGND VPWR VPWR net1980 sky130_fd_sc_hd__dlygate4sd3_1
X_14248_ clknet_leaf_258_clk _02877_ VGND VGND VPWR VPWR data_array.data1\[12\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_78_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14179_ clknet_leaf_238_clk _02808_ VGND VGND VPWR VPWR data_array.data0\[2\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_125_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout809 net810 VGND VGND VPWR VPWR net809 sky130_fd_sc_hd__clkbuf_4
XFILLER_113_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08740_ net764 net2960 net463 VGND VGND VPWR VPWR _00499_ sky130_fd_sc_hd__mux2_1
XFILLER_79_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1007 tag_array.tag1\[12\]\[11\] VGND VGND VPWR VPWR net2658 sky130_fd_sc_hd__dlygate4sd3_1
X_05952_ data_array.rdata1\[40\] net1657 net843 VGND VGND VPWR VPWR _03429_ sky130_fd_sc_hd__a21o_1
Xhold1018 tag_array.tag0\[8\]\[16\] VGND VGND VPWR VPWR net2669 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1029 data_array.data0\[3\]\[37\] VGND VGND VPWR VPWR net2680 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1380 net1382 VGND VGND VPWR VPWR net1380 sky130_fd_sc_hd__clkbuf_2
X_08671_ net740 net4221 net501 VGND VGND VPWR VPWR _00430_ sky130_fd_sc_hd__mux2_1
Xfanout1391 net1392 VGND VGND VPWR VPWR net1391 sky130_fd_sc_hd__clkbuf_4
X_05883_ data_array.rdata1\[17\] net829 net838 VGND VGND VPWR VPWR _03383_ sky130_fd_sc_hd__a21o_1
X_07622_ data_array.data1\[12\]\[16\] net1353 net1259 data_array.data1\[15\]\[16\]
+ _04846_ VGND VGND VPWR VPWR _04847_ sky130_fd_sc_hd__a221o_1
XFILLER_66_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07553_ data_array.data1\[5\]\[10\] net1604 net1508 data_array.data1\[6\]\[10\] VGND
+ VGND VPWR VPWR _04784_ sky130_fd_sc_hd__a22o_1
XFILLER_179_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06504_ net1172 _03825_ _03829_ net1221 VGND VGND VPWR VPWR _03831_ sky130_fd_sc_hd__a22o_1
XFILLER_179_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07484_ _04720_ _04721_ VGND VGND VPWR VPWR _00097_ sky130_fd_sc_hd__or2_1
XFILLER_146_1064 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_3377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09223_ net789 net2932 net645 VGND VGND VPWR VPWR _00977_ sky130_fd_sc_hd__mux2_1
XFILLER_166_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_3388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06435_ tag_array.tag0\[1\]\[22\] net1562 net1466 tag_array.tag0\[2\]\[22\] VGND
+ VGND VPWR VPWR _03768_ sky130_fd_sc_hd__a22o_1
XFILLER_107_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09154_ net924 net3202 net566 VGND VGND VPWR VPWR _00908_ sky130_fd_sc_hd__mux2_1
X_06366_ tag_array.tag0\[4\]\[16\] net1408 net1314 tag_array.tag0\[7\]\[16\] _03704_
+ VGND VGND VPWR VPWR _03705_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_118_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_650 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08105_ data_array.data1\[13\]\[60\] net1604 net1508 data_array.data1\[14\]\[60\]
+ VGND VGND VPWR VPWR _05286_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_135_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09085_ net946 net4318 net410 VGND VGND VPWR VPWR _00839_ sky130_fd_sc_hd__mux2_1
X_06297_ tag_array.tag0\[13\]\[10\] net1596 net1500 tag_array.tag0\[14\]\[10\] VGND
+ VGND VPWR VPWR _03642_ sky130_fd_sc_hd__a22o_1
XFILLER_174_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08036_ data_array.data1\[8\]\[54\] net1355 net1261 data_array.data1\[11\]\[54\]
+ _05222_ VGND VGND VPWR VPWR _05223_ sky130_fd_sc_hd__a221o_1
XFILLER_107_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput90 cpu_wdata[60] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_1
XFILLER_116_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold830 data_array.data0\[1\]\[29\] VGND VGND VPWR VPWR net2481 sky130_fd_sc_hd__dlygate4sd3_1
Xhold841 tag_array.tag1\[11\]\[0\] VGND VGND VPWR VPWR net2492 sky130_fd_sc_hd__dlygate4sd3_1
Xhold852 tag_array.tag0\[9\]\[22\] VGND VGND VPWR VPWR net2503 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold863 data_array.data0\[2\]\[31\] VGND VGND VPWR VPWR net2514 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_153_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold874 tag_array.tag0\[13\]\[13\] VGND VGND VPWR VPWR net2525 sky130_fd_sc_hd__dlygate4sd3_1
Xhold885 data_array.data1\[3\]\[63\] VGND VGND VPWR VPWR net2536 sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 tag_array.tag1\[1\]\[4\] VGND VGND VPWR VPWR net2547 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_1076 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09987_ net880 net4200 net374 VGND VGND VPWR VPWR _01736_ sky130_fd_sc_hd__mux2_1
Xhold2220 data_array.data0\[12\]\[17\] VGND VGND VPWR VPWR net3871 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2231 data_array.data1\[9\]\[37\] VGND VGND VPWR VPWR net3882 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2242 tag_array.tag1\[15\]\[20\] VGND VGND VPWR VPWR net3893 sky130_fd_sc_hd__dlygate4sd3_1
X_08938_ net1012 net2543 net432 VGND VGND VPWR VPWR _00694_ sky130_fd_sc_hd__mux2_1
Xhold2253 tag_array.tag0\[14\]\[11\] VGND VGND VPWR VPWR net3904 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2264 data_array.data1\[3\]\[3\] VGND VGND VPWR VPWR net3915 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1530 data_array.data1\[12\]\[51\] VGND VGND VPWR VPWR net3181 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2275 data_array.data0\[5\]\[63\] VGND VGND VPWR VPWR net3926 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1541 data_array.data1\[3\]\[13\] VGND VGND VPWR VPWR net3192 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2286 tag_array.tag0\[6\]\[24\] VGND VGND VPWR VPWR net3937 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2297 tag_array.tag1\[6\]\[16\] VGND VGND VPWR VPWR net3948 sky130_fd_sc_hd__dlygate4sd3_1
X_08869_ net1028 net2562 net440 VGND VGND VPWR VPWR _00626_ sky130_fd_sc_hd__mux2_1
Xhold1552 tag_array.tag1\[10\]\[21\] VGND VGND VPWR VPWR net3203 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1563 data_array.data0\[8\]\[4\] VGND VGND VPWR VPWR net3214 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1574 tag_array.tag1\[15\]\[4\] VGND VGND VPWR VPWR net3225 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1585 data_array.data1\[11\]\[26\] VGND VGND VPWR VPWR net3236 sky130_fd_sc_hd__dlygate4sd3_1
X_10900_ net886 net3624 net515 VGND VGND VPWR VPWR _02645_ sky130_fd_sc_hd__mux2_1
XFILLER_85_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11880_ clknet_leaf_48_clk _00688_ VGND VGND VPWR VPWR data_array.data0\[5\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1596 tag_array.tag1\[3\]\[12\] VGND VGND VPWR VPWR net3247 sky130_fd_sc_hd__dlygate4sd3_1
X_10831_ net2163 net906 net502 VGND VGND VPWR VPWR _02576_ sky130_fd_sc_hd__mux2_1
XFILLER_16_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13550_ clknet_leaf_78_clk _02179_ VGND VGND VPWR VPWR data_array.data1\[0\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_41_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10762_ net924 net4011 net490 VGND VGND VPWR VPWR _02507_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12501_ clknet_leaf_5_clk _01195_ VGND VGND VPWR VPWR data_array.data1\[9\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
X_13481_ clknet_leaf_154_clk _02111_ VGND VGND VPWR VPWR tag_array.tag0\[15\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_10693_ net2790 net944 net478 VGND VGND VPWR VPWR _02438_ sky130_fd_sc_hd__mux2_1
XFILLER_13_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12432_ clknet_leaf_25_clk _01126_ VGND VGND VPWR VPWR data_array.data0\[14\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12363_ clknet_leaf_14_clk _00039_ VGND VGND VPWR VPWR data_array.rdata0\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14102_ clknet_leaf_49_clk _02731_ VGND VGND VPWR VPWR data_array.data0\[1\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_154_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11314_ net1039 net4004 net796 VGND VGND VPWR VPWR _03057_ sky130_fd_sc_hd__mux2_1
XFILLER_180_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12294_ clknet_leaf_167_clk _01052_ VGND VGND VPWR VPWR tag_array.tag1\[12\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14033_ clknet_leaf_58_clk _02662_ VGND VGND VPWR VPWR data_array.data1\[6\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_11245_ net1050 net2549 net681 VGND VGND VPWR VPWR _02988_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11176_ net1070 net3669 net658 VGND VGND VPWR VPWR _02919_ sky130_fd_sc_hd__mux2_1
XFILLER_164_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10127_ net1037 net3580 net363 VGND VGND VPWR VPWR _01875_ sky130_fd_sc_hd__mux2_1
XFILLER_48_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10058_ net793 net3046 net600 VGND VGND VPWR VPWR _01807_ sky130_fd_sc_hd__mux2_1
XFILLER_169_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13817_ clknet_leaf_55_clk _02446_ VGND VGND VPWR VPWR data_array.data1\[2\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_995 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13748_ clknet_leaf_83_clk _02377_ VGND VGND VPWR VPWR data_array.data1\[1\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13679_ clknet_leaf_240_clk _02308_ VGND VGND VPWR VPWR data_array.data1\[15\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_14_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06220_ tag_array.tag0\[13\]\[3\] net1564 net1468 tag_array.tag0\[14\]\[3\] VGND
+ VGND VPWR VPWR _03572_ sky130_fd_sc_hd__a22o_1
XFILLER_31_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06151_ net27 net26 VGND VGND VPWR VPWR _03508_ sky130_fd_sc_hd__and2b_4
XTAP_TAPCELL_ROW_152_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold104 data_array.data0\[2\]\[40\] VGND VGND VPWR VPWR net1755 sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 data_array.data1\[0\]\[13\] VGND VGND VPWR VPWR net1766 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold126 tag_array.tag1\[1\]\[21\] VGND VGND VPWR VPWR net1777 sky130_fd_sc_hd__dlygate4sd3_1
X_06082_ fsm.tag_out0\[23\] net1121 _03504_ VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_113_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold137 data_array.data1\[2\]\[63\] VGND VGND VPWR VPWR net1788 sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 data_array.data1\[2\]\[62\] VGND VGND VPWR VPWR net1799 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_99_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09910_ net769 net4584 net602 VGND VGND VPWR VPWR _01660_ sky130_fd_sc_hd__mux2_1
Xhold159 tag_array.dirty1\[0\] VGND VGND VPWR VPWR net1810 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout606 net608 VGND VGND VPWR VPWR net606 sky130_fd_sc_hd__buf_4
X_09841_ net1105 net4245 net378 VGND VGND VPWR VPWR _01591_ sky130_fd_sc_hd__mux2_1
Xfanout617 _05571_ VGND VGND VPWR VPWR net617 sky130_fd_sc_hd__buf_2
Xfanout628 net629 VGND VGND VPWR VPWR net628 sky130_fd_sc_hd__buf_4
XFILLER_58_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_615 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout639 net644 VGND VGND VPWR VPWR net639 sky130_fd_sc_hd__clkbuf_8
XFILLER_140_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09772_ net3985 net701 net672 VGND VGND VPWR VPWR _01524_ sky130_fd_sc_hd__mux2_1
X_06984_ data_array.data0\[12\]\[22\] net1341 net1247 data_array.data0\[15\]\[22\]
+ _04266_ VGND VGND VPWR VPWR _04267_ sky130_fd_sc_hd__a221o_1
X_08723_ net1758 net730 net474 VGND VGND VPWR VPWR _00482_ sky130_fd_sc_hd__mux2_1
X_05935_ net126 net1151 _03416_ _03417_ VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__a22o_1
XFILLER_67_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08654_ net1892 net706 net511 VGND VGND VPWR VPWR _00413_ sky130_fd_sc_hd__mux2_1
X_05866_ net101 net1156 _03371_ _03370_ VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_159_3417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07605_ _04830_ _04831_ VGND VGND VPWR VPWR _00069_ sky130_fd_sc_hd__or2_1
XFILLER_81_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08585_ net782 net2968 net530 VGND VGND VPWR VPWR _00344_ sky130_fd_sc_hd__mux2_1
XFILLER_54_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_05797_ _03309_ _03310_ _03311_ _03313_ VGND VGND VPWR VPWR _03314_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_176_3742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07536_ data_array.data1\[0\]\[8\] net1345 net1251 data_array.data1\[3\]\[8\] _04768_
+ VGND VGND VPWR VPWR _04769_ sky130_fd_sc_hd__a221o_1
XFILLER_169_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07467_ data_array.data1\[9\]\[2\] net1526 net1430 data_array.data1\[10\]\[2\] VGND
+ VGND VPWR VPWR _04706_ sky130_fd_sc_hd__a22o_1
XFILLER_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09206_ net755 net3118 net631 VGND VGND VPWR VPWR _00960_ sky130_fd_sc_hd__mux2_1
X_06418_ tag_array.tag0\[13\]\[21\] net1600 net1504 tag_array.tag0\[14\]\[21\] VGND
+ VGND VPWR VPWR _03752_ sky130_fd_sc_hd__a22o_1
X_07398_ data_array.data0\[8\]\[60\] net1414 net1320 data_array.data0\[11\]\[60\]
+ _04642_ VGND VGND VPWR VPWR _04643_ sky130_fd_sc_hd__a221o_1
XFILLER_10_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_1012 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09137_ net995 net4188 net573 VGND VGND VPWR VPWR _00891_ sky130_fd_sc_hd__mux2_1
X_06349_ net1625 _03683_ _03687_ net1199 VGND VGND VPWR VPWR _03690_ sky130_fd_sc_hd__a22o_1
XFILLER_136_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09068_ net1012 net3392 net414 VGND VGND VPWR VPWR _00822_ sky130_fd_sc_hd__mux2_1
XFILLER_118_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08019_ data_array.data1\[1\]\[52\] net1545 net1449 data_array.data1\[2\]\[52\] VGND
+ VGND VPWR VPWR _05208_ sky130_fd_sc_hd__a22o_1
Xhold660 data_array.data0\[14\]\[62\] VGND VGND VPWR VPWR net2311 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_420 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold671 data_array.data0\[8\]\[16\] VGND VGND VPWR VPWR net2322 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_5_13__f_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_5_13__leaf_clk sky130_fd_sc_hd__clkbuf_16
Xhold682 data_array.data0\[2\]\[63\] VGND VGND VPWR VPWR net2333 sky130_fd_sc_hd__dlygate4sd3_1
X_11030_ net3713 net880 net340 VGND VGND VPWR VPWR _02774_ sky130_fd_sc_hd__mux2_1
Xhold693 tag_array.tag1\[4\]\[5\] VGND VGND VPWR VPWR net2344 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2050 tag_array.tag1\[5\]\[17\] VGND VGND VPWR VPWR net3701 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2061 data_array.data0\[11\]\[54\] VGND VGND VPWR VPWR net3712 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2072 data_array.data1\[6\]\[50\] VGND VGND VPWR VPWR net3723 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_40_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2083 tag_array.tag0\[7\]\[15\] VGND VGND VPWR VPWR net3734 sky130_fd_sc_hd__dlygate4sd3_1
X_12981_ clknet_leaf_156_clk _01675_ VGND VGND VPWR VPWR tag_array.tag0\[4\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_134_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2094 tag_array.tag1\[13\]\[23\] VGND VGND VPWR VPWR net3745 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1360 tag_array.tag0\[8\]\[0\] VGND VGND VPWR VPWR net3011 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1371 tag_array.tag0\[14\]\[17\] VGND VGND VPWR VPWR net3022 sky130_fd_sc_hd__dlygate4sd3_1
X_11932_ clknet_leaf_270_clk _00740_ VGND VGND VPWR VPWR data_array.data0\[4\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1382 data_array.data1\[0\]\[54\] VGND VGND VPWR VPWR net3033 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1393 data_array.data0\[10\]\[46\] VGND VGND VPWR VPWR net3044 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11863_ clknet_leaf_262_clk _00671_ VGND VGND VPWR VPWR data_array.data0\[5\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_150_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10814_ net1917 net974 net503 VGND VGND VPWR VPWR _02559_ sky130_fd_sc_hd__mux2_1
X_13602_ clknet_leaf_230_clk _02231_ VGND VGND VPWR VPWR data_array.data0\[9\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_0_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11794_ clknet_leaf_115_clk _00602_ VGND VGND VPWR VPWR data_array.data0\[8\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13533_ clknet_leaf_69_clk _02162_ VGND VGND VPWR VPWR data_array.data1\[0\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10745_ net994 net4353 net496 VGND VGND VPWR VPWR _02490_ sky130_fd_sc_hd__mux2_1
XFILLER_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13464_ clknet_leaf_168_clk _02094_ VGND VGND VPWR VPWR tag_array.tag0\[1\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_97_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10676_ net3290 net1015 net485 VGND VGND VPWR VPWR _02421_ sky130_fd_sc_hd__mux2_1
XFILLER_127_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12415_ clknet_leaf_72_clk _01109_ VGND VGND VPWR VPWR data_array.data0\[14\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
X_13395_ clknet_leaf_70_clk _02025_ VGND VGND VPWR VPWR data_array.data1\[8\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_58_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12346_ clknet_leaf_14_clk _00020_ VGND VGND VPWR VPWR data_array.rdata0\[28\] sky130_fd_sc_hd__dfxtp_1
Xoutput209 net209 VGND VGND VPWR VPWR cpu_rdata[4] sky130_fd_sc_hd__buf_6
XFILLER_182_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12277_ clknet_leaf_127_clk _01035_ VGND VGND VPWR VPWR tag_array.tag1\[13\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_126_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14016_ clknet_leaf_13_clk _02645_ VGND VGND VPWR VPWR data_array.data1\[5\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
X_11228_ net863 net2540 net658 VGND VGND VPWR VPWR _02971_ sky130_fd_sc_hd__mux2_1
XFILLER_96_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11159_ net883 net3076 net542 VGND VGND VPWR VPWR _02902_ sky130_fd_sc_hd__mux2_1
XFILLER_96_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05720_ net14 fsm.tag_out1\[14\] VGND VGND VPWR VPWR _03237_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_19_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05651_ fsm.tag_out0\[0\] net30 VGND VGND VPWR VPWR _03168_ sky130_fd_sc_hd__and2b_1
XFILLER_63_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08370_ net124 net59 net1639 VGND VGND VPWR VPWR _05483_ sky130_fd_sc_hd__mux2_1
XFILLER_51_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07321_ data_array.data0\[8\]\[53\] net1334 net1240 data_array.data0\[11\]\[53\]
+ _04572_ VGND VGND VPWR VPWR _04573_ sky130_fd_sc_hd__a221o_1
XFILLER_17_1026 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07252_ net1168 _04505_ _04509_ net1216 VGND VGND VPWR VPWR _04511_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_171_3650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06203_ tag_array.tag0\[12\]\[1\] net1402 net1308 tag_array.tag0\[15\]\[1\] _03556_
+ VGND VGND VPWR VPWR _03557_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_30_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07183_ data_array.data0\[1\]\[40\] net1603 net1507 data_array.data0\[2\]\[40\] VGND
+ VGND VPWR VPWR _04448_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_30_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_132_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06134_ data_array.rdata0\[49\] net1140 net1114 data_array.rdata1\[49\] VGND VGND
+ VPWR VPWR net306 sky130_fd_sc_hd__a22o_1
XFILLER_172_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06065_ net1161 net15 fsm.tag_out1\[15\] net1132 VGND VGND VPWR VPWR _03496_ sky130_fd_sc_hd__a22o_1
Xfanout403 net409 VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__buf_4
XFILLER_132_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout414 net415 VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__buf_4
Xfanout425 _05610_ VGND VGND VPWR VPWR net425 sky130_fd_sc_hd__clkbuf_8
Xfanout436 net437 VGND VGND VPWR VPWR net436 sky130_fd_sc_hd__buf_4
XFILLER_98_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout447 net448 VGND VGND VPWR VPWR net447 sky130_fd_sc_hd__buf_4
X_09824_ net913 net3126 net391 VGND VGND VPWR VPWR _01575_ sky130_fd_sc_hd__mux2_1
Xfanout458 net459 VGND VGND VPWR VPWR net458 sky130_fd_sc_hd__buf_4
Xfanout469 net470 VGND VGND VPWR VPWR net469 sky130_fd_sc_hd__buf_4
XFILLER_101_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_12 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06967_ _04250_ _04251_ VGND VGND VPWR VPWR _00012_ sky130_fd_sc_hd__or2_1
X_09755_ net2357 net766 net664 VGND VGND VPWR VPWR _01507_ sky130_fd_sc_hd__mux2_1
XFILLER_100_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08706_ net2296 net700 net488 VGND VGND VPWR VPWR _00465_ sky130_fd_sc_hd__mux2_1
X_05918_ data_array.rdata0\[29\] net1658 net1148 VGND VGND VPWR VPWR _03406_ sky130_fd_sc_hd__o21a_1
X_09686_ net744 net3585 net605 VGND VGND VPWR VPWR _01438_ sky130_fd_sc_hd__mux2_1
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06898_ data_array.data0\[0\]\[14\] net1378 net1284 data_array.data0\[3\]\[14\] _04188_
+ VGND VGND VPWR VPWR _04189_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_169_Left_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08637_ net2237 net774 net505 VGND VGND VPWR VPWR _00396_ sky130_fd_sc_hd__mux2_1
X_05849_ data_array.rdata0\[6\] net846 net1142 VGND VGND VPWR VPWR _03360_ sky130_fd_sc_hd__o21a_1
XFILLER_70_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08568_ net811 _05577_ VGND VGND VPWR VPWR _05599_ sky130_fd_sc_hd__nand2_2
XFILLER_168_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07519_ data_array.data1\[8\]\[7\] net1398 net1304 data_array.data1\[11\]\[7\] _04752_
+ VGND VGND VPWR VPWR _04753_ sky130_fd_sc_hd__a221o_1
XFILLER_11_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08499_ net1722 net618 VGND VGND VPWR VPWR _00295_ sky130_fd_sc_hd__nand2b_1
X_10530_ net1086 net3938 net453 VGND VGND VPWR VPWR _02275_ sky130_fd_sc_hd__mux2_1
XFILLER_183_704 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10461_ net1103 net2615 net346 VGND VGND VPWR VPWR _02206_ sky130_fd_sc_hd__mux2_1
XFILLER_164_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12200_ clknet_leaf_145_clk _00153_ VGND VGND VPWR VPWR fsm.tag_out0\[7\] sky130_fd_sc_hd__dfxtp_2
XPHY_EDGE_ROW_178_Left_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13180_ clknet_leaf_253_clk _00072_ VGND VGND VPWR VPWR data_array.rdata1\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10392_ net3014 net1086 net661 VGND VGND VPWR VPWR _02138_ sky130_fd_sc_hd__mux2_1
XFILLER_135_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12131_ clknet_leaf_145_clk _00939_ VGND VGND VPWR VPWR tag_array.tag0\[12\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_53_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12062_ clknet_leaf_19_clk _00870_ VGND VGND VPWR VPWR data_array.data1\[14\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold490 data_array.data0\[4\]\[35\] VGND VGND VPWR VPWR net2141 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_151_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11013_ net1854 net948 net343 VGND VGND VPWR VPWR _02757_ sky130_fd_sc_hd__mux2_1
XFILLER_49_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout970 net971 VGND VGND VPWR VPWR net970 sky130_fd_sc_hd__clkbuf_2
Xfanout981 _05484_ VGND VGND VPWR VPWR net981 sky130_fd_sc_hd__buf_1
Xfanout992 _05478_ VGND VGND VPWR VPWR net992 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12964_ clknet_leaf_177_clk _01658_ VGND VGND VPWR VPWR tag_array.tag0\[4\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_79_1031 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1190 data_array.data0\[7\]\[53\] VGND VGND VPWR VPWR net2841 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11915_ clknet_leaf_2_clk _00723_ VGND VGND VPWR VPWR data_array.data0\[5\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12895_ clknet_leaf_225_clk _01589_ VGND VGND VPWR VPWR data_array.data0\[12\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1078 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11846_ clknet_leaf_40_clk _00654_ VGND VGND VPWR VPWR data_array.data0\[7\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11777_ clknet_leaf_46_clk _00585_ VGND VGND VPWR VPWR data_array.data0\[8\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
X_13516_ clknet_leaf_200_clk _02145_ VGND VGND VPWR VPWR data_array.data1\[0\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_10728_ net1062 net4098 net498 VGND VGND VPWR VPWR _02473_ sky130_fd_sc_hd__mux2_1
X_14496_ clknet_leaf_161_clk _03119_ VGND VGND VPWR VPWR tag_array.dirty0\[14\] sky130_fd_sc_hd__dfxtp_1
X_10659_ net2577 net1083 net485 VGND VGND VPWR VPWR _02404_ sky130_fd_sc_hd__mux2_1
X_13447_ clknet_leaf_176_clk _02077_ VGND VGND VPWR VPWR tag_array.tag0\[1\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload13 clknet_5_28__leaf_clk VGND VGND VPWR VPWR clkload13/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload24 clknet_leaf_263_clk VGND VGND VPWR VPWR clkload24/Y sky130_fd_sc_hd__clkinv_8
Xclkload35 clknet_leaf_16_clk VGND VGND VPWR VPWR clkload35/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload46 clknet_leaf_256_clk VGND VGND VPWR VPWR clkload46/Y sky130_fd_sc_hd__bufinv_16
XFILLER_6_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13378_ clknet_leaf_108_clk _02008_ VGND VGND VPWR VPWR tag_array.tag0\[2\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload57 clknet_leaf_255_clk VGND VGND VPWR VPWR clkload57/Y sky130_fd_sc_hd__inv_6
XFILLER_170_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload68 clknet_leaf_233_clk VGND VGND VPWR VPWR clkload68/Y sky130_fd_sc_hd__inv_12
Xclkload79 clknet_leaf_51_clk VGND VGND VPWR VPWR clkload79/Y sky130_fd_sc_hd__inv_6
X_12329_ clknet_leaf_49_clk _00002_ VGND VGND VPWR VPWR data_array.rdata0\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_48_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2808 tag_array.tag0\[1\]\[22\] VGND VGND VPWR VPWR net4459 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2819 data_array.data0\[13\]\[0\] VGND VGND VPWR VPWR net4470 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07870_ data_array.data1\[9\]\[39\] net1538 net1442 data_array.data1\[10\]\[39\]
+ VGND VGND VPWR VPWR _05072_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_147_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06821_ data_array.data0\[4\]\[7\] net1411 net1317 data_array.data0\[7\]\[7\] _04118_
+ VGND VGND VPWR VPWR _04119_ sky130_fd_sc_hd__a221o_1
XFILLER_28_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09540_ net768 net3657 net618 VGND VGND VPWR VPWR _01293_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_108_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06752_ data_array.data0\[9\]\[1\] net1523 net1427 data_array.data0\[10\]\[1\] VGND
+ VGND VPWR VPWR _04056_ sky130_fd_sc_hd__a22o_1
XFILLER_37_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05703_ net30 net1655 VGND VGND VPWR VPWR _03220_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_125_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09471_ net742 net4204 net654 VGND VGND VPWR VPWR _01224_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_125_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06683_ tag_array.tag1\[8\]\[20\] net1368 net1274 tag_array.tag1\[11\]\[20\] _03992_
+ VGND VGND VPWR VPWR _03993_ sky130_fd_sc_hd__a221o_1
XFILLER_93_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08422_ net1127 _05517_ VGND VGND VPWR VPWR _05518_ sky130_fd_sc_hd__and2_1
X_05634_ net4625 _03151_ _03152_ VGND VGND VPWR VPWR _00188_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_121_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08353_ net1123 _05471_ VGND VGND VPWR VPWR _05472_ sky130_fd_sc_hd__and2_1
X_07304_ data_array.data0\[1\]\[51\] net1522 net1426 data_array.data0\[2\]\[51\] VGND
+ VGND VPWR VPWR _04558_ sky130_fd_sc_hd__a22o_1
XFILLER_20_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_178_Right_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08284_ net1128 _05425_ VGND VGND VPWR VPWR _05426_ sky130_fd_sc_hd__and2_1
Xclkload7 clknet_5_14__leaf_clk VGND VGND VPWR VPWR clkload7/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_149_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07235_ data_array.data0\[0\]\[45\] net1344 net1250 data_array.data0\[3\]\[45\] _04494_
+ VGND VGND VPWR VPWR _04495_ sky130_fd_sc_hd__a221o_1
XFILLER_166_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07166_ data_array.data0\[9\]\[39\] net1541 net1445 data_array.data0\[10\]\[39\]
+ VGND VGND VPWR VPWR _04432_ sky130_fd_sc_hd__a22o_1
XFILLER_133_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06117_ data_array.rdata0\[32\] net1134 net1113 data_array.rdata1\[32\] VGND VGND
+ VPWR VPWR net288 sky130_fd_sc_hd__a22o_1
X_07097_ net1188 _04363_ _04367_ net1614 VGND VGND VPWR VPWR _04370_ sky130_fd_sc_hd__a22o_1
XFILLER_132_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06048_ fsm.tag_out0\[6\] net1120 _03487_ VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__a21o_1
XFILLER_59_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1209 net1211 VGND VGND VPWR VPWR net1209 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_184_3885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_184_3896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09807_ net983 net3003 net386 VGND VGND VPWR VPWR _01558_ sky130_fd_sc_hd__mux2_1
X_07999_ net1616 _05183_ _05187_ net1190 VGND VGND VPWR VPWR _05190_ sky130_fd_sc_hd__a22o_1
XFILLER_86_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09738_ net734 net4093 net679 VGND VGND VPWR VPWR _01490_ sky130_fd_sc_hd__mux2_1
XFILLER_74_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09669_ net712 net3602 net612 VGND VGND VPWR VPWR _01421_ sky130_fd_sc_hd__mux2_1
X_11700_ clknet_leaf_136_clk _00508_ VGND VGND VPWR VPWR tag_array.tag1\[15\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_12680_ clknet_leaf_110_clk _01374_ VGND VGND VPWR VPWR data_array.data0\[15\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11631_ clknet_leaf_196_clk _00439_ VGND VGND VPWR VPWR tag_array.tag1\[3\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_46_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_145_Right_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11562_ clknet_leaf_191_clk _00370_ VGND VGND VPWR VPWR tag_array.tag1\[5\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_14350_ clknet_leaf_174_clk _02973_ VGND VGND VPWR VPWR data_array.data1\[10\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10513_ net894 net3434 net346 VGND VGND VPWR VPWR _02258_ sky130_fd_sc_hd__mux2_1
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13301_ clknet_leaf_111_clk _01931_ VGND VGND VPWR VPWR data_array.data0\[10\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_14281_ clknet_leaf_265_clk _02910_ VGND VGND VPWR VPWR data_array.data1\[11\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_11493_ clknet_leaf_153_clk _00302_ VGND VGND VPWR VPWR tag_array.valid0\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_183_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_567 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13232_ clknet_leaf_204_clk _01862_ VGND VGND VPWR VPWR data_array.data0\[11\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_21_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10444_ net1983 net878 net665 VGND VGND VPWR VPWR _02190_ sky130_fd_sc_hd__mux2_1
XFILLER_108_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13163_ clknet_leaf_185_clk _00064_ VGND VGND VPWR VPWR data_array.rdata1\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10375_ net699 net2120 net539 VGND VGND VPWR VPWR _02122_ sky130_fd_sc_hd__mux2_1
XFILLER_136_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12114_ clknet_leaf_119_clk _00922_ VGND VGND VPWR VPWR data_array.data1\[14\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
X_13094_ clknet_leaf_28_clk _01788_ VGND VGND VPWR VPWR data_array.data1\[13\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_152_998 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12045_ clknet_leaf_14_clk _00853_ VGND VGND VPWR VPWR data_array.data0\[6\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_49_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13996_ clknet_leaf_82_clk _02625_ VGND VGND VPWR VPWR data_array.data1\[5\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_46_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_142_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12947_ clknet_leaf_1_clk _01641_ VGND VGND VPWR VPWR data_array.data0\[13\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_66_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12878_ clknet_leaf_23_clk _01572_ VGND VGND VPWR VPWR data_array.data0\[12\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_103_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_367 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11829_ clknet_leaf_34_clk _00637_ VGND VGND VPWR VPWR data_array.data0\[7\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_112_Right_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14479_ clknet_leaf_204_clk _03102_ VGND VGND VPWR VPWR data_array.data1\[7\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload102 clknet_leaf_37_clk VGND VGND VPWR VPWR clkload102/Y sky130_fd_sc_hd__inv_6
Xclkload113 clknet_leaf_96_clk VGND VGND VPWR VPWR clkload113/Y sky130_fd_sc_hd__inv_6
XFILLER_162_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07020_ net1188 _04293_ _04297_ net1614 VGND VGND VPWR VPWR _04300_ sky130_fd_sc_hd__a22o_1
Xclkload124 clknet_leaf_79_clk VGND VGND VPWR VPWR clkload124/Y sky130_fd_sc_hd__inv_8
Xclkload135 clknet_leaf_217_clk VGND VGND VPWR VPWR clkload135/Y sky130_fd_sc_hd__inv_8
Xclkload146 clknet_leaf_211_clk VGND VGND VPWR VPWR clkload146/Y sky130_fd_sc_hd__bufinv_16
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload157 clknet_leaf_170_clk VGND VGND VPWR VPWR clkload157/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_155_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload168 clknet_leaf_206_clk VGND VGND VPWR VPWR clkload168/X sky130_fd_sc_hd__clkbuf_4
Xclkload179 clknet_leaf_179_clk VGND VGND VPWR VPWR clkload179/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_149_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08971_ net882 net2553 net429 VGND VGND VPWR VPWR _00727_ sky130_fd_sc_hd__mux2_1
XFILLER_88_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_166_3560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2605 data_array.data0\[7\]\[11\] VGND VGND VPWR VPWR net4256 sky130_fd_sc_hd__dlygate4sd3_1
X_07922_ net1628 _05113_ _05117_ net1202 VGND VGND VPWR VPWR _05120_ sky130_fd_sc_hd__a22o_1
Xhold2616 data_array.data0\[13\]\[29\] VGND VGND VPWR VPWR net4267 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2627 tag_array.tag1\[5\]\[21\] VGND VGND VPWR VPWR net4278 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2638 tag_array.tag0\[8\]\[15\] VGND VGND VPWR VPWR net4289 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2649 tag_array.tag1\[9\]\[23\] VGND VGND VPWR VPWR net4300 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1904 data_array.data0\[13\]\[44\] VGND VGND VPWR VPWR net3555 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_127_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1915 data_array.data0\[13\]\[25\] VGND VGND VPWR VPWR net3566 sky130_fd_sc_hd__dlygate4sd3_1
X_07853_ data_array.data1\[12\]\[37\] net1353 net1259 data_array.data1\[15\]\[37\]
+ _05056_ VGND VGND VPWR VPWR _05057_ sky130_fd_sc_hd__a221o_1
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1926 data_array.data1\[0\]\[37\] VGND VGND VPWR VPWR net3577 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_162_3468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1937 tag_array.tag0\[7\]\[17\] VGND VGND VPWR VPWR net3588 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_162_3479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1948 tag_array.tag1\[11\]\[16\] VGND VGND VPWR VPWR net3599 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06804_ data_array.data0\[8\]\[6\] net1332 net1238 data_array.data0\[11\]\[6\] _04102_
+ VGND VGND VPWR VPWR _04103_ sky130_fd_sc_hd__a221o_1
Xhold1959 tag_array.tag0\[15\]\[3\] VGND VGND VPWR VPWR net3610 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07784_ data_array.data1\[5\]\[31\] net1574 net1478 data_array.data1\[6\]\[31\] VGND
+ VGND VPWR VPWR _04994_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06735_ net1172 _04035_ _04039_ net1221 VGND VGND VPWR VPWR _04041_ sky130_fd_sc_hd__a22o_1
X_09523_ net737 net3268 net621 VGND VGND VPWR VPWR _01276_ sky130_fd_sc_hd__mux2_1
XFILLER_36_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09454_ net819 net4090 _05568_ VGND VGND VPWR VPWR _01207_ sky130_fd_sc_hd__mux2_1
X_06666_ tag_array.tag1\[5\]\[18\] net1562 net1466 tag_array.tag1\[6\]\[18\] VGND
+ VGND VPWR VPWR _03978_ sky130_fd_sc_hd__a22o_1
XFILLER_101_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05617_ net10 VGND VGND VPWR VPWR _03139_ sky130_fd_sc_hd__inv_2
X_08405_ net2254 net936 net692 VGND VGND VPWR VPWR _00264_ sky130_fd_sc_hd__mux2_1
X_09385_ net861 net2311 net409 VGND VGND VPWR VPWR _01138_ sky130_fd_sc_hd__mux2_1
X_06597_ tag_array.tag1\[4\]\[12\] net1401 net1307 tag_array.tag1\[7\]\[12\] _03914_
+ VGND VGND VPWR VPWR _03915_ sky130_fd_sc_hd__a221o_1
X_08336_ net2837 net1028 net693 VGND VGND VPWR VPWR _00241_ sky130_fd_sc_hd__mux2_1
XFILLER_184_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08267_ fsm.tag_out1\[24\] net816 net808 fsm.tag_out0\[24\] _05412_ VGND VGND VPWR
+ VPWR _05413_ sky130_fd_sc_hd__a221o_1
XFILLER_137_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_140_clk clknet_5_31__leaf_clk VGND VGND VPWR VPWR clknet_leaf_140_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_124_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07218_ net1628 _04473_ _04477_ net1202 VGND VGND VPWR VPWR _04480_ sky130_fd_sc_hd__a22o_1
XFILLER_137_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_717 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08198_ fsm.tag_out1\[1\] net816 net808 fsm.tag_out0\[1\] _05366_ VGND VGND VPWR
+ VPWR _05367_ sky130_fd_sc_hd__a221o_1
XFILLER_106_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07149_ data_array.data0\[12\]\[37\] net1356 net1262 data_array.data0\[15\]\[37\]
+ _04416_ VGND VGND VPWR VPWR _04417_ sky130_fd_sc_hd__a221o_1
XFILLER_118_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_762 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10160_ net905 net3418 net362 VGND VGND VPWR VPWR _01908_ sky130_fd_sc_hd__mux2_1
XFILLER_10_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1006 net1007 VGND VGND VPWR VPWR net1006 sky130_fd_sc_hd__clkbuf_2
XFILLER_117_1039 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1017 _05466_ VGND VGND VPWR VPWR net1017 sky130_fd_sc_hd__buf_1
X_10091_ net1816 net760 net643 VGND VGND VPWR VPWR _01840_ sky130_fd_sc_hd__mux2_1
Xfanout1028 _05460_ VGND VGND VPWR VPWR net1028 sky130_fd_sc_hd__clkbuf_2
Xfanout1039 _05456_ VGND VGND VPWR VPWR net1039 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_76_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13850_ clknet_leaf_18_clk _02479_ VGND VGND VPWR VPWR data_array.data1\[3\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12801_ clknet_leaf_103_clk _01495_ VGND VGND VPWR VPWR tag_array.tag1\[10\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10993_ net2859 net1028 net343 VGND VGND VPWR VPWR _02737_ sky130_fd_sc_hd__mux2_1
X_13781_ clknet_leaf_200_clk _02410_ VGND VGND VPWR VPWR data_array.data1\[2\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_48_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_643 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12732_ clknet_leaf_105_clk _01426_ VGND VGND VPWR VPWR tag_array.tag0\[5\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_805 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ clknet_leaf_20_clk _01357_ VGND VGND VPWR VPWR data_array.data0\[15\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_26_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14402_ clknet_leaf_213_clk _03025_ VGND VGND VPWR VPWR data_array.data1\[10\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_169_873 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11614_ clknet_leaf_135_clk _00422_ VGND VGND VPWR VPWR tag_array.tag1\[3\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_61_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12594_ clknet_leaf_166_clk _01288_ VGND VGND VPWR VPWR tag_array.tag0\[0\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_169_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_85_Right_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14333_ clknet_leaf_5_clk _02962_ VGND VGND VPWR VPWR data_array.data1\[11\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
X_11545_ clknet_leaf_33_clk _00353_ VGND VGND VPWR VPWR tag_array.tag1\[6\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_131_clk clknet_5_30__leaf_clk VGND VGND VPWR VPWR clknet_leaf_131_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_51_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14264_ clknet_leaf_75_clk _02893_ VGND VGND VPWR VPWR data_array.data1\[12\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
X_11476_ clknet_leaf_175_clk _00286_ VGND VGND VPWR VPWR tag_array.valid1\[0\] sky130_fd_sc_hd__dfxtp_1
X_10427_ net1946 net944 net661 VGND VGND VPWR VPWR _02173_ sky130_fd_sc_hd__mux2_1
X_13215_ clknet_leaf_212_clk _00111_ VGND VGND VPWR VPWR data_array.rdata1\[52\] sky130_fd_sc_hd__dfxtp_1
X_14195_ clknet_leaf_49_clk _02824_ VGND VGND VPWR VPWR data_array.data0\[2\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_151_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10358_ net768 net4259 net540 VGND VGND VPWR VPWR _02105_ sky130_fd_sc_hd__mux2_1
X_13146_ clknet_leaf_137_clk _01840_ VGND VGND VPWR VPWR tag_array.tag1\[8\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_151_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13077_ clknet_leaf_30_clk _01771_ VGND VGND VPWR VPWR data_array.data1\[13\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10289_ net1757 net1005 net634 VGND VGND VPWR VPWR _02036_ sky130_fd_sc_hd__mux2_1
XFILLER_140_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_94_Right_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12028_ clknet_leaf_89_clk _00836_ VGND VGND VPWR VPWR data_array.data0\[6\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout1540 net1542 VGND VGND VPWR VPWR net1540 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_144_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1551 net1554 VGND VGND VPWR VPWR net1551 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_144_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_198_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_198_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_39_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1562 net1563 VGND VGND VPWR VPWR net1562 sky130_fd_sc_hd__clkbuf_4
XFILLER_78_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1573 net1591 VGND VGND VPWR VPWR net1573 sky130_fd_sc_hd__clkbuf_2
Xfanout1584 net1591 VGND VGND VPWR VPWR net1584 sky130_fd_sc_hd__clkbuf_4
XFILLER_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1595 net1596 VGND VGND VPWR VPWR net1595 sky130_fd_sc_hd__clkbuf_4
XFILLER_25_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13979_ clknet_leaf_66_clk _02608_ VGND VGND VPWR VPWR data_array.data1\[5\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_06520_ tag_array.tag1\[0\]\[5\] net1420 net1326 tag_array.tag1\[3\]\[5\] _03844_
+ VGND VGND VPWR VPWR _03845_ sky130_fd_sc_hd__a221o_1
XFILLER_179_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06451_ tag_array.tag0\[9\]\[24\] net1565 net1469 tag_array.tag0\[10\]\[24\] VGND
+ VGND VPWR VPWR _03782_ sky130_fd_sc_hd__a22o_1
XFILLER_15_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09170_ net863 net2215 net576 VGND VGND VPWR VPWR _00924_ sky130_fd_sc_hd__mux2_1
XFILLER_166_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06382_ net1208 _03713_ _03717_ net1634 VGND VGND VPWR VPWR _03720_ sky130_fd_sc_hd__a22o_1
XFILLER_21_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08121_ net1219 _05295_ _05299_ net1171 VGND VGND VPWR VPWR _05301_ sky130_fd_sc_hd__a22o_1
XFILLER_119_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_122_clk clknet_5_27__leaf_clk VGND VGND VPWR VPWR clknet_leaf_122_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_179_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08052_ data_array.data1\[5\]\[55\] net1534 net1438 data_array.data1\[6\]\[55\] VGND
+ VGND VPWR VPWR _05238_ sky130_fd_sc_hd__a22o_1
XFILLER_135_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07003_ data_array.data0\[5\]\[24\] net1578 net1482 data_array.data0\[6\]\[24\] VGND
+ VGND VPWR VPWR _04284_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_116_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2402 tag_array.tag0\[2\]\[2\] VGND VGND VPWR VPWR net4053 sky130_fd_sc_hd__dlygate4sd3_1
Xinput109 mem_rdata[19] VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__clkbuf_1
Xhold2413 data_array.data1\[14\]\[41\] VGND VGND VPWR VPWR net4064 sky130_fd_sc_hd__dlygate4sd3_1
X_08954_ net948 net2696 net432 VGND VGND VPWR VPWR _00710_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_181_3833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2424 data_array.data0\[13\]\[56\] VGND VGND VPWR VPWR net4075 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_181_3844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2435 data_array.data1\[6\]\[49\] VGND VGND VPWR VPWR net4086 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2446 data_array.data1\[10\]\[62\] VGND VGND VPWR VPWR net4097 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_5_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1701 data_array.data1\[15\]\[11\] VGND VGND VPWR VPWR net3352 sky130_fd_sc_hd__dlygate4sd3_1
X_07905_ data_array.data1\[5\]\[42\] net1586 net1490 data_array.data1\[6\]\[42\] VGND
+ VGND VPWR VPWR _05104_ sky130_fd_sc_hd__a22o_1
Xhold1712 data_array.data0\[5\]\[1\] VGND VGND VPWR VPWR net3363 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2457 tag_array.tag1\[15\]\[0\] VGND VGND VPWR VPWR net4108 sky130_fd_sc_hd__dlygate4sd3_1
X_08885_ net964 net3688 net440 VGND VGND VPWR VPWR _00642_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_189_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_189_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_56_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1723 tag_array.tag0\[8\]\[2\] VGND VGND VPWR VPWR net3374 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2468 data_array.data0\[13\]\[43\] VGND VGND VPWR VPWR net4119 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1734 data_array.data1\[12\]\[28\] VGND VGND VPWR VPWR net3385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2479 data_array.data0\[12\]\[51\] VGND VGND VPWR VPWR net4130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1745 tag_array.tag0\[1\]\[8\] VGND VGND VPWR VPWR net3396 sky130_fd_sc_hd__dlygate4sd3_1
X_07836_ _05040_ _05041_ VGND VGND VPWR VPWR _00092_ sky130_fd_sc_hd__or2_1
Xhold1756 tag_array.tag0\[11\]\[1\] VGND VGND VPWR VPWR net3407 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1767 data_array.data0\[11\]\[51\] VGND VGND VPWR VPWR net3418 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1778 data_array.data1\[7\]\[50\] VGND VGND VPWR VPWR net3429 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1789 lru_array.lru_mem\[12\] VGND VGND VPWR VPWR net3440 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_16_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_12 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_34 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07767_ data_array.data1\[4\]\[29\] net1382 net1288 data_array.data1\[7\]\[29\] _04978_
+ VGND VGND VPWR VPWR _04979_ sky130_fd_sc_hd__a221o_1
X_09506_ net704 net2747 _05565_ VGND VGND VPWR VPWR _01259_ sky130_fd_sc_hd__mux2_1
X_06718_ tag_array.tag1\[4\]\[23\] net1419 net1325 tag_array.tag1\[7\]\[23\] _04024_
+ VGND VGND VPWR VPWR _04025_ sky130_fd_sc_hd__a221o_1
X_07698_ data_array.data1\[9\]\[23\] net1553 net1457 data_array.data1\[10\]\[23\]
+ VGND VGND VPWR VPWR _04916_ sky130_fd_sc_hd__a22o_1
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_179_3795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09437_ net919 net4168 net586 VGND VGND VPWR VPWR _01190_ sky130_fd_sc_hd__mux2_1
X_06649_ tag_array.tag1\[13\]\[17\] net1609 net1513 tag_array.tag1\[14\]\[17\] VGND
+ VGND VPWR VPWR _03962_ sky130_fd_sc_hd__a22o_1
XFILLER_169_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09368_ net929 net4618 net403 VGND VGND VPWR VPWR _01121_ sky130_fd_sc_hd__mux2_1
XFILLER_162_1070 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08319_ net105 net40 net1640 VGND VGND VPWR VPWR _05449_ sky130_fd_sc_hd__mux2_1
X_09299_ net783 net3012 net544 VGND VGND VPWR VPWR _01053_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_113_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_113_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_166_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_60 net1495 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_71 _00084_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_82 net1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11330_ net974 net3862 net796 VGND VGND VPWR VPWR _03073_ sky130_fd_sc_hd__mux2_1
XANTENNA_93 net1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11261_ net984 net4390 net680 VGND VGND VPWR VPWR _03004_ sky130_fd_sc_hd__mux2_1
XFILLER_21_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10212_ net957 net4599 net359 VGND VGND VPWR VPWR _01959_ sky130_fd_sc_hd__mux2_1
X_13000_ clknet_leaf_63_clk _01694_ VGND VGND VPWR VPWR data_array.data0\[3\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_11192_ net1005 net3236 net649 VGND VGND VPWR VPWR _02935_ sky130_fd_sc_hd__mux2_1
X_10143_ net973 net3175 net362 VGND VGND VPWR VPWR _01891_ sky130_fd_sc_hd__mux2_1
X_10074_ net726 net3435 net601 VGND VGND VPWR VPWR _01823_ sky130_fd_sc_hd__mux2_1
X_13902_ clknet_leaf_269_clk _02531_ VGND VGND VPWR VPWR data_array.data1\[4\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_85_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13833_ clknet_leaf_266_clk _02462_ VGND VGND VPWR VPWR data_array.data1\[3\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13764_ clknet_leaf_115_clk _02393_ VGND VGND VPWR VPWR data_array.data1\[1\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
X_10976_ net1928 net1096 net342 VGND VGND VPWR VPWR _02720_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_100_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12715_ clknet_leaf_144_clk _01409_ VGND VGND VPWR VPWR tag_array.tag0\[7\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_13695_ clknet_leaf_20_clk _02324_ VGND VGND VPWR VPWR data_array.data1\[15\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_80_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12646_ clknet_leaf_31_clk _01340_ VGND VGND VPWR VPWR data_array.data0\[15\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_104_clk clknet_5_24__leaf_clk VGND VGND VPWR VPWR clknet_leaf_104_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_156_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12577_ clknet_leaf_158_clk _01271_ VGND VGND VPWR VPWR tag_array.tag0\[10\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_172_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14316_ clknet_leaf_118_clk _02945_ VGND VGND VPWR VPWR data_array.data1\[11\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_172_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11528_ clknet_leaf_174_clk _00336_ VGND VGND VPWR VPWR tag_array.valid1\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_117_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_846 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold308 data_array.data1\[1\]\[6\] VGND VGND VPWR VPWR net1959 sky130_fd_sc_hd__dlygate4sd3_1
Xhold319 data_array.data0\[2\]\[28\] VGND VGND VPWR VPWR net1970 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_78_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14247_ clknet_leaf_37_clk _02876_ VGND VGND VPWR VPWR data_array.data1\[12\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_171_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11459_ clknet_leaf_40_clk _00269_ VGND VGND VPWR VPWR data_array.data0\[0\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_78_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_123_Left_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14178_ clknet_leaf_246_clk _02807_ VGND VGND VPWR VPWR data_array.data0\[2\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_124_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13129_ clknet_leaf_157_clk _01823_ VGND VGND VPWR VPWR tag_array.tag0\[3\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_05951_ data_array.rdata0\[40\] net1659 net1149 VGND VGND VPWR VPWR _03428_ sky130_fd_sc_hd__o21a_1
Xhold1008 data_array.data1\[12\]\[2\] VGND VGND VPWR VPWR net2659 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1019 data_array.data1\[11\]\[3\] VGND VGND VPWR VPWR net2670 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_223 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1370 net1376 VGND VGND VPWR VPWR net1370 sky130_fd_sc_hd__clkbuf_2
X_08670_ net742 net3247 net501 VGND VGND VPWR VPWR _00429_ sky130_fd_sc_hd__mux2_1
X_05882_ data_array.rdata0\[17\] net847 net1142 VGND VGND VPWR VPWR _03382_ sky130_fd_sc_hd__o21a_1
Xfanout1381 net1382 VGND VGND VPWR VPWR net1381 sky130_fd_sc_hd__clkbuf_4
XFILLER_27_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1392 net1400 VGND VGND VPWR VPWR net1392 sky130_fd_sc_hd__clkbuf_2
XFILLER_26_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07621_ data_array.data1\[13\]\[16\] net1544 net1448 data_array.data1\[14\]\[16\]
+ VGND VGND VPWR VPWR _04846_ sky130_fd_sc_hd__a22o_1
XFILLER_26_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_132_Left_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07552_ data_array.data1\[8\]\[10\] net1414 net1320 data_array.data1\[11\]\[10\]
+ _04782_ VGND VGND VPWR VPWR _04783_ sky130_fd_sc_hd__a221o_1
X_06503_ net1623 _03823_ _03827_ net1197 VGND VGND VPWR VPWR _03830_ sky130_fd_sc_hd__a22o_1
XFILLER_50_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07483_ net1177 _04715_ _04719_ net1225 VGND VGND VPWR VPWR _04721_ sky130_fd_sc_hd__a22o_1
XFILLER_146_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_3378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06434_ tag_array.tag0\[12\]\[22\] net1374 net1280 tag_array.tag0\[15\]\[22\] _03766_
+ VGND VGND VPWR VPWR _03767_ sky130_fd_sc_hd__a221o_1
X_09222_ net793 net3276 net646 VGND VGND VPWR VPWR _00976_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_157_3389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09153_ net930 net4225 net568 VGND VGND VPWR VPWR _00907_ sky130_fd_sc_hd__mux2_1
X_06365_ tag_array.tag0\[5\]\[16\] net1600 net1504 tag_array.tag0\[6\]\[16\] VGND
+ VGND VPWR VPWR _03704_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_118_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08104_ data_array.data1\[4\]\[60\] net1414 net1320 data_array.data1\[7\]\[60\] _05284_
+ VGND VGND VPWR VPWR _05285_ sky130_fd_sc_hd__a221o_1
XFILLER_163_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09084_ net948 net3302 net416 VGND VGND VPWR VPWR _00838_ sky130_fd_sc_hd__mux2_1
X_06296_ _03640_ _03641_ VGND VGND VPWR VPWR _00155_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_135_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_141_Left_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08035_ data_array.data1\[9\]\[54\] net1544 net1448 data_array.data1\[10\]\[54\]
+ VGND VGND VPWR VPWR _05222_ sky130_fd_sc_hd__a22o_1
XFILLER_162_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold820 data_array.data0\[5\]\[9\] VGND VGND VPWR VPWR net2471 sky130_fd_sc_hd__dlygate4sd3_1
Xinput80 cpu_wdata[51] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_1
XFILLER_116_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput91 cpu_wdata[61] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_1
Xhold831 tag_array.tag1\[2\]\[2\] VGND VGND VPWR VPWR net2482 sky130_fd_sc_hd__dlygate4sd3_1
Xhold842 data_array.data1\[15\]\[60\] VGND VGND VPWR VPWR net2493 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold853 tag_array.tag1\[1\]\[17\] VGND VGND VPWR VPWR net2504 sky130_fd_sc_hd__dlygate4sd3_1
Xhold864 data_array.data0\[2\]\[39\] VGND VGND VPWR VPWR net2515 sky130_fd_sc_hd__dlygate4sd3_1
Xhold875 tag_array.tag0\[6\]\[3\] VGND VGND VPWR VPWR net2526 sky130_fd_sc_hd__dlygate4sd3_1
Xhold886 tag_array.tag1\[3\]\[10\] VGND VGND VPWR VPWR net2537 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold897 tag_array.tag1\[9\]\[22\] VGND VGND VPWR VPWR net2548 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09986_ net884 net4480 net371 VGND VGND VPWR VPWR _01735_ sky130_fd_sc_hd__mux2_1
Xhold2210 tag_array.tag0\[9\]\[4\] VGND VGND VPWR VPWR net3861 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2221 tag_array.tag1\[11\]\[13\] VGND VGND VPWR VPWR net3872 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2232 data_array.data0\[10\]\[59\] VGND VGND VPWR VPWR net3883 sky130_fd_sc_hd__dlygate4sd3_1
X_08937_ net1018 net3675 net429 VGND VGND VPWR VPWR _00693_ sky130_fd_sc_hd__mux2_1
Xhold2243 tag_array.tag0\[0\]\[3\] VGND VGND VPWR VPWR net3894 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2254 data_array.data1\[7\]\[39\] VGND VGND VPWR VPWR net3905 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2265 tag_array.tag0\[5\]\[24\] VGND VGND VPWR VPWR net3916 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1520 data_array.data1\[0\]\[28\] VGND VGND VPWR VPWR net3171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2276 data_array.data0\[7\]\[46\] VGND VGND VPWR VPWR net3927 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1531 tag_array.tag1\[4\]\[14\] VGND VGND VPWR VPWR net3182 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2287 data_array.data1\[15\]\[6\] VGND VGND VPWR VPWR net3938 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1542 data_array.data0\[5\]\[53\] VGND VGND VPWR VPWR net3193 sky130_fd_sc_hd__dlygate4sd3_1
X_08868_ net1032 net4180 net438 VGND VGND VPWR VPWR _00625_ sky130_fd_sc_hd__mux2_1
Xhold1553 data_array.data1\[11\]\[43\] VGND VGND VPWR VPWR net3204 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2298 tag_array.tag1\[13\]\[6\] VGND VGND VPWR VPWR net3949 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_150_Left_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1564 data_array.data1\[4\]\[16\] VGND VGND VPWR VPWR net3215 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1575 data_array.data0\[5\]\[8\] VGND VGND VPWR VPWR net3226 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_83_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1586 data_array.data0\[9\]\[62\] VGND VGND VPWR VPWR net3237 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_28_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07819_ data_array.data1\[9\]\[34\] net1532 net1436 data_array.data1\[10\]\[34\]
+ VGND VGND VPWR VPWR _05026_ sky130_fd_sc_hd__a22o_1
XFILLER_72_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1597 data_array.data0\[9\]\[30\] VGND VGND VPWR VPWR net3248 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08799_ net1761 net1049 net447 VGND VGND VPWR VPWR _00557_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10830_ net1900 net908 net504 VGND VGND VPWR VPWR _02575_ sky130_fd_sc_hd__mux2_1
XFILLER_44_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10761_ net930 net3119 net492 VGND VGND VPWR VPWR _02506_ sky130_fd_sc_hd__mux2_1
XFILLER_16_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12500_ clknet_leaf_212_clk _01194_ VGND VGND VPWR VPWR data_array.data1\[9\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10692_ net1919 net950 net487 VGND VGND VPWR VPWR _02437_ sky130_fd_sc_hd__mux2_1
X_13480_ clknet_leaf_163_clk _02110_ VGND VGND VPWR VPWR tag_array.tag0\[15\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_12431_ clknet_leaf_53_clk _01125_ VGND VGND VPWR VPWR data_array.data0\[14\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12362_ clknet_leaf_81_clk _00038_ VGND VGND VPWR VPWR data_array.rdata0\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_154_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14101_ clknet_leaf_225_clk _02730_ VGND VGND VPWR VPWR data_array.data0\[1\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_153_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11313_ net1040 net3131 net795 VGND VGND VPWR VPWR _03056_ sky130_fd_sc_hd__mux2_1
X_12293_ clknet_leaf_96_clk _01051_ VGND VGND VPWR VPWR tag_array.tag1\[12\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_181_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14032_ clknet_leaf_28_clk _02661_ VGND VGND VPWR VPWR data_array.data1\[6\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_11244_ net1055 net2529 net680 VGND VGND VPWR VPWR _02987_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11175_ net1075 net4002 net656 VGND VGND VPWR VPWR _02918_ sky130_fd_sc_hd__mux2_1
X_10126_ net1043 net2591 net362 VGND VGND VPWR VPWR _01874_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_73_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10057_ net859 net3773 net558 VGND VGND VPWR VPWR _01806_ sky130_fd_sc_hd__mux2_1
XFILLER_57_82 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1076 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13816_ clknet_leaf_75_clk _02445_ VGND VGND VPWR VPWR data_array.data1\[2\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
X_13747_ clknet_leaf_36_clk _02376_ VGND VGND VPWR VPWR data_array.data1\[1\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_139_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10959_ net906 net4218 net526 VGND VGND VPWR VPWR _02704_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_139_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13678_ clknet_leaf_77_clk _02307_ VGND VGND VPWR VPWR data_array.data1\[15\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_14_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12629_ clknet_leaf_45_clk _01323_ VGND VGND VPWR VPWR data_array.data0\[15\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06150_ net28 net29 VGND VGND VPWR VPWR _03507_ sky130_fd_sc_hd__nand2b_1
XFILLER_89_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold105 tag_array.tag1\[0\]\[22\] VGND VGND VPWR VPWR net1756 sky130_fd_sc_hd__dlygate4sd3_1
X_06081_ net1164 net24 fsm.tag_out1\[23\] net1133 VGND VGND VPWR VPWR _03504_ sky130_fd_sc_hd__a22o_1
XFILLER_172_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_113_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold116 data_array.data0\[8\]\[49\] VGND VGND VPWR VPWR net1767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 data_array.data0\[8\]\[7\] VGND VGND VPWR VPWR net1778 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 tag_array.tag1\[0\]\[5\] VGND VGND VPWR VPWR net1789 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold149 data_array.data1\[8\]\[45\] VGND VGND VPWR VPWR net1800 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_125_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09840_ net1109 net4470 net381 VGND VGND VPWR VPWR _01590_ sky130_fd_sc_hd__mux2_1
Xfanout607 net608 VGND VGND VPWR VPWR net607 sky130_fd_sc_hd__buf_2
Xfanout618 net620 VGND VGND VPWR VPWR net618 sky130_fd_sc_hd__buf_4
Xfanout629 _05563_ VGND VGND VPWR VPWR net629 sky130_fd_sc_hd__buf_4
XFILLER_86_627 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09771_ net1756 net702 net665 VGND VGND VPWR VPWR _01523_ sky130_fd_sc_hd__mux2_1
X_06983_ data_array.data0\[13\]\[22\] net1532 net1436 data_array.data0\[14\]\[22\]
+ VGND VGND VPWR VPWR _04266_ sky130_fd_sc_hd__a22o_1
XFILLER_86_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08722_ net2750 net735 net470 VGND VGND VPWR VPWR _00481_ sky130_fd_sc_hd__mux2_1
X_05934_ data_array.rdata1\[34\] net829 net838 VGND VGND VPWR VPWR _03417_ sky130_fd_sc_hd__a21o_1
X_08653_ net2339 net711 net503 VGND VGND VPWR VPWR _00412_ sky130_fd_sc_hd__mux2_1
X_05865_ data_array.rdata1\[11\] net833 net842 VGND VGND VPWR VPWR _03371_ sky130_fd_sc_hd__a21o_1
XFILLER_96_1048 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_3418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07604_ net1176 _04825_ _04829_ net1225 VGND VGND VPWR VPWR _04831_ sky130_fd_sc_hd__a22o_1
X_08584_ net786 net2510 net537 VGND VGND VPWR VPWR _00343_ sky130_fd_sc_hd__mux2_1
X_05796_ _03280_ _03282_ _03312_ VGND VGND VPWR VPWR _03313_ sky130_fd_sc_hd__or3_1
XFILLER_81_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_176_3743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07535_ data_array.data1\[1\]\[8\] net1535 net1439 data_array.data1\[2\]\[8\] VGND
+ VGND VPWR VPWR _04768_ sky130_fd_sc_hd__a22o_1
XFILLER_35_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07466_ data_array.data1\[4\]\[2\] net1336 net1242 data_array.data1\[7\]\[2\] _04704_
+ VGND VGND VPWR VPWR _04705_ sky130_fd_sc_hd__a221o_1
X_06417_ _03750_ _03751_ VGND VGND VPWR VPWR _00143_ sky130_fd_sc_hd__or2_1
X_09205_ net759 net2563 net632 VGND VGND VPWR VPWR _00959_ sky130_fd_sc_hd__mux2_1
X_07397_ data_array.data0\[9\]\[60\] net1604 net1508 data_array.data0\[10\]\[60\]
+ VGND VGND VPWR VPWR _04642_ sky130_fd_sc_hd__a22o_1
XFILLER_33_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06348_ tag_array.tag0\[0\]\[14\] net1368 net1274 tag_array.tag0\[3\]\[14\] _03688_
+ VGND VGND VPWR VPWR _03689_ sky130_fd_sc_hd__a221o_1
X_09136_ net999 net3170 net569 VGND VGND VPWR VPWR _00890_ sky130_fd_sc_hd__mux2_1
XFILLER_176_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09067_ net1018 net3474 net413 VGND VGND VPWR VPWR _00821_ sky130_fd_sc_hd__mux2_1
XFILLER_120_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06279_ tag_array.tag0\[13\]\[8\] net1599 net1503 tag_array.tag0\[14\]\[8\] VGND
+ VGND VPWR VPWR _03626_ sky130_fd_sc_hd__a22o_1
X_08018_ data_array.data1\[8\]\[52\] net1354 net1260 data_array.data1\[11\]\[52\]
+ _05206_ VGND VGND VPWR VPWR _05207_ sky130_fd_sc_hd__a221o_1
Xhold650 data_array.data1\[3\]\[19\] VGND VGND VPWR VPWR net2301 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_151_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_326 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold661 tag_array.tag0\[14\]\[15\] VGND VGND VPWR VPWR net2312 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold672 data_array.data0\[5\]\[35\] VGND VGND VPWR VPWR net2323 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold683 data_array.data0\[7\]\[2\] VGND VGND VPWR VPWR net2334 sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 data_array.data0\[0\]\[28\] VGND VGND VPWR VPWR net2345 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_34_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09969_ net955 net3932 net374 VGND VGND VPWR VPWR _01718_ sky130_fd_sc_hd__mux2_1
Xhold2040 tag_array.tag1\[15\]\[8\] VGND VGND VPWR VPWR net3691 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2051 tag_array.tag1\[6\]\[23\] VGND VGND VPWR VPWR net3702 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2062 data_array.data0\[1\]\[57\] VGND VGND VPWR VPWR net3713 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12980_ clknet_leaf_169_clk _01674_ VGND VGND VPWR VPWR tag_array.tag0\[4\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2073 data_array.data0\[4\]\[40\] VGND VGND VPWR VPWR net3724 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_182_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2084 data_array.data0\[10\]\[56\] VGND VGND VPWR VPWR net3735 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1350 tag_array.tag1\[4\]\[8\] VGND VGND VPWR VPWR net3001 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2095 data_array.data1\[13\]\[0\] VGND VGND VPWR VPWR net3746 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1047 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1361 tag_array.tag1\[12\]\[2\] VGND VGND VPWR VPWR net3012 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1372 tag_array.tag1\[12\]\[17\] VGND VGND VPWR VPWR net3023 sky130_fd_sc_hd__dlygate4sd3_1
X_11931_ clknet_leaf_210_clk _00739_ VGND VGND VPWR VPWR data_array.data0\[4\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1383 tag_array.tag1\[14\]\[20\] VGND VGND VPWR VPWR net3034 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1394 tag_array.tag0\[7\]\[14\] VGND VGND VPWR VPWR net3045 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11862_ clknet_leaf_230_clk _00670_ VGND VGND VPWR VPWR data_array.data0\[5\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_13601_ clknet_leaf_242_clk _02230_ VGND VGND VPWR VPWR data_array.data0\[9\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_10813_ net2181 net978 net509 VGND VGND VPWR VPWR _02558_ sky130_fd_sc_hd__mux2_1
XFILLER_14_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11793_ clknet_leaf_54_clk _00601_ VGND VGND VPWR VPWR data_array.data0\[8\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
X_13532_ clknet_leaf_40_clk _02161_ VGND VGND VPWR VPWR data_array.data1\[0\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_10744_ net997 net4605 net492 VGND VGND VPWR VPWR _02489_ sky130_fd_sc_hd__mux2_1
XFILLER_159_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13463_ clknet_leaf_102_clk _02093_ VGND VGND VPWR VPWR tag_array.tag0\[1\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_10675_ net2201 net1016 net481 VGND VGND VPWR VPWR _02420_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_97_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12414_ clknet_leaf_261_clk _01108_ VGND VGND VPWR VPWR data_array.data0\[14\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
X_13394_ clknet_leaf_42_clk _02024_ VGND VGND VPWR VPWR data_array.data1\[8\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_58_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12345_ clknet_leaf_215_clk _00019_ VGND VGND VPWR VPWR data_array.rdata0\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_126_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12276_ clknet_leaf_137_clk _01034_ VGND VGND VPWR VPWR tag_array.tag1\[13\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_14015_ clknet_leaf_17_clk _02644_ VGND VGND VPWR VPWR data_array.data1\[5\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
X_11227_ net864 net4041 net652 VGND VGND VPWR VPWR _02970_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11158_ net887 net2522 net543 VGND VGND VPWR VPWR _02901_ sky130_fd_sc_hd__mux2_1
XFILLER_110_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10109_ net1108 net3943 net365 VGND VGND VPWR VPWR _01857_ sky130_fd_sc_hd__mux2_1
X_11089_ net2107 net904 net328 VGND VGND VPWR VPWR _02832_ sky130_fd_sc_hd__mux2_1
XFILLER_64_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_159_Right_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05650_ net20 fsm.tag_out0\[20\] VGND VGND VPWR VPWR _03167_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_19_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07320_ data_array.data0\[9\]\[53\] net1531 net1435 data_array.data0\[10\]\[53\]
+ VGND VGND VPWR VPWR _04572_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_154_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1038 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07251_ net1618 _04503_ _04507_ net1192 VGND VGND VPWR VPWR _04510_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_171_3640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_171_3651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06202_ tag_array.tag0\[13\]\[1\] net1559 net1463 tag_array.tag0\[14\]\[1\] VGND
+ VGND VPWR VPWR _03556_ sky130_fd_sc_hd__a22o_1
X_07182_ data_array.data0\[8\]\[40\] net1415 net1321 data_array.data0\[11\]\[40\]
+ _04446_ VGND VGND VPWR VPWR _04447_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_30_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06133_ data_array.rdata0\[48\] net1141 net1116 data_array.rdata1\[48\] VGND VGND
+ VPWR VPWR net305 sky130_fd_sc_hd__a22o_1
XFILLER_145_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06064_ fsm.tag_out0\[14\] net1120 _03495_ VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__a21o_1
XFILLER_117_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout404 net405 VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__clkbuf_8
XFILLER_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout415 net417 VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__buf_4
Xfanout426 net433 VGND VGND VPWR VPWR net426 sky130_fd_sc_hd__clkbuf_8
XFILLER_86_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout437 net441 VGND VGND VPWR VPWR net437 sky130_fd_sc_hd__buf_4
X_09823_ net916 net2978 net391 VGND VGND VPWR VPWR _01574_ sky130_fd_sc_hd__mux2_1
Xfanout448 net449 VGND VGND VPWR VPWR net448 sky130_fd_sc_hd__clkbuf_8
Xfanout459 _05604_ VGND VGND VPWR VPWR net459 sky130_fd_sc_hd__clkbuf_4
XFILLER_140_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09754_ net1789 net772 net671 VGND VGND VPWR VPWR _01506_ sky130_fd_sc_hd__mux2_1
X_06966_ net1184 _04245_ _04249_ net1232 VGND VGND VPWR VPWR _04251_ sky130_fd_sc_hd__a22o_1
XFILLER_104_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08705_ net1747 net702 net482 VGND VGND VPWR VPWR _00464_ sky130_fd_sc_hd__mux2_1
X_05917_ net119 net1151 _03404_ _03405_ VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__a22o_1
X_09685_ net748 net3686 net605 VGND VGND VPWR VPWR _01437_ sky130_fd_sc_hd__mux2_1
X_06897_ data_array.data0\[1\]\[14\] net1567 net1471 data_array.data0\[2\]\[14\] VGND
+ VGND VPWR VPWR _04188_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_93_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_93_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_126_Right_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08636_ net3364 net778 net506 VGND VGND VPWR VPWR _00395_ sky130_fd_sc_hd__mux2_1
X_05848_ net154 net1153 _03358_ _03359_ VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__a22o_1
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08567_ net811 _05574_ net1695 VGND VGND VPWR VPWR _00334_ sky130_fd_sc_hd__a21o_1
X_05779_ fsm.tag_out1\[4\] net3 VGND VGND VPWR VPWR _03296_ sky130_fd_sc_hd__and2b_1
XFILLER_70_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07518_ data_array.data1\[9\]\[7\] net1589 net1493 data_array.data1\[10\]\[7\] VGND
+ VGND VPWR VPWR _04752_ sky130_fd_sc_hd__a22o_1
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08498_ net821 net812 net854 _05416_ VGND VGND VPWR VPWR _05569_ sky130_fd_sc_hd__or4b_1
X_07449_ net1199 _04683_ _04687_ net1625 VGND VGND VPWR VPWR _04690_ sky130_fd_sc_hd__a22o_1
XFILLER_183_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xwire827 _03333_ VGND VGND VPWR VPWR net827 sky130_fd_sc_hd__clkbuf_2
XFILLER_182_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10460_ net1105 net4601 net344 VGND VGND VPWR VPWR _02205_ sky130_fd_sc_hd__mux2_1
X_09119_ net1066 net3153 net573 VGND VGND VPWR VPWR _00873_ sky130_fd_sc_hd__mux2_1
XFILLER_136_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10391_ net2419 net1090 net664 VGND VGND VPWR VPWR _02137_ sky130_fd_sc_hd__mux2_1
XFILLER_136_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_92_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12130_ clknet_leaf_154_clk _00938_ VGND VGND VPWR VPWR tag_array.tag0\[12\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_92_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_53_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12061_ clknet_leaf_82_clk _00869_ VGND VGND VPWR VPWR data_array.data1\[14\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_53_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold480 data_array.data0\[8\]\[12\] VGND VGND VPWR VPWR net2131 sky130_fd_sc_hd__dlygate4sd3_1
Xhold491 tag_array.tag1\[1\]\[13\] VGND VGND VPWR VPWR net2142 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11012_ net2468 net954 net340 VGND VGND VPWR VPWR _02756_ sky130_fd_sc_hd__mux2_1
XFILLER_145_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout960 net963 VGND VGND VPWR VPWR net960 sky130_fd_sc_hd__clkbuf_2
XFILLER_77_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout971 _05490_ VGND VGND VPWR VPWR net971 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout982 _05484_ VGND VGND VPWR VPWR net982 sky130_fd_sc_hd__clkbuf_2
Xfanout993 _05478_ VGND VGND VPWR VPWR net993 sky130_fd_sc_hd__buf_1
XFILLER_18_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_5_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12963_ clknet_leaf_177_clk _01657_ VGND VGND VPWR VPWR tag_array.tag0\[4\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_92_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_84_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_84_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_79_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1180 tag_array.tag0\[8\]\[17\] VGND VGND VPWR VPWR net2831 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1191 data_array.data0\[12\]\[53\] VGND VGND VPWR VPWR net2842 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11914_ clknet_leaf_213_clk _00722_ VGND VGND VPWR VPWR data_array.data0\[5\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
X_12894_ clknet_leaf_110_clk _01588_ VGND VGND VPWR VPWR data_array.data0\[12\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11845_ clknet_leaf_91_clk _00653_ VGND VGND VPWR VPWR data_array.data0\[7\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11776_ clknet_leaf_93_clk _00584_ VGND VGND VPWR VPWR data_array.data0\[8\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
X_13515_ clknet_leaf_85_clk _02144_ VGND VGND VPWR VPWR data_array.data1\[0\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_10727_ net1067 net4079 net496 VGND VGND VPWR VPWR _02472_ sky130_fd_sc_hd__mux2_1
X_14495_ clknet_leaf_176_clk _03118_ VGND VGND VPWR VPWR lru_array.lru_mem\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_70_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13446_ clknet_leaf_168_clk _02076_ VGND VGND VPWR VPWR tag_array.tag0\[1\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_10658_ net3308 net1086 net478 VGND VGND VPWR VPWR _02403_ sky130_fd_sc_hd__mux2_1
XFILLER_139_470 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload14 clknet_5_30__leaf_clk VGND VGND VPWR VPWR clkload14/Y sky130_fd_sc_hd__inv_6
Xclkload25 clknet_leaf_264_clk VGND VGND VPWR VPWR clkload25/Y sky130_fd_sc_hd__inv_8
Xclkload36 clknet_leaf_17_clk VGND VGND VPWR VPWR clkload36/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_86_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload47 clknet_leaf_257_clk VGND VGND VPWR VPWR clkload47/Y sky130_fd_sc_hd__clkinv_2
X_13377_ clknet_leaf_191_clk _02007_ VGND VGND VPWR VPWR tag_array.tag0\[2\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_10589_ net2630 net1104 net466 VGND VGND VPWR VPWR _02334_ sky130_fd_sc_hd__mux2_1
Xclkload58 clknet_leaf_24_clk VGND VGND VPWR VPWR clkload58/X sky130_fd_sc_hd__clkbuf_8
XFILLER_6_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload69 clknet_leaf_235_clk VGND VGND VPWR VPWR clkload69/Y sky130_fd_sc_hd__inv_8
XFILLER_126_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12328_ clknet_leaf_119_clk _00001_ VGND VGND VPWR VPWR data_array.rdata0\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_115_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12259_ clknet_leaf_136_clk _01017_ VGND VGND VPWR VPWR tag_array.tag1\[14\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2809 data_array.data1\[3\]\[53\] VGND VGND VPWR VPWR net4460 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_95_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_147_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06820_ data_array.data0\[5\]\[7\] net1601 net1505 data_array.data0\[6\]\[7\] VGND
+ VGND VPWR VPWR _04118_ sky130_fd_sc_hd__a22o_1
XFILLER_96_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1020 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_416 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06751_ data_array.data0\[0\]\[1\] net1333 net1239 data_array.data0\[3\]\[1\] _04054_
+ VGND VGND VPWR VPWR _04055_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_108_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_75_clk clknet_5_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_75_clk sky130_fd_sc_hd__clkbuf_8
X_05702_ _03187_ _03188_ _03218_ VGND VGND VPWR VPWR _03219_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_125_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06682_ tag_array.tag1\[9\]\[20\] net1558 net1462 tag_array.tag1\[10\]\[20\] VGND
+ VGND VPWR VPWR _03992_ sky130_fd_sc_hd__a22o_1
X_09470_ net747 net3899 net655 VGND VGND VPWR VPWR _01223_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_125_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08421_ net142 net77 net1641 VGND VGND VPWR VPWR _05517_ sky130_fd_sc_hd__mux2_1
X_05633_ net1158 net327 net1649 VGND VGND VPWR VPWR _03152_ sky130_fd_sc_hd__mux2_1
XFILLER_24_549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08352_ net117 net52 net1639 VGND VGND VPWR VPWR _05471_ sky130_fd_sc_hd__mux2_1
X_07303_ data_array.data0\[8\]\[51\] net1332 net1238 data_array.data0\[11\]\[51\]
+ _04556_ VGND VGND VPWR VPWR _04557_ sky130_fd_sc_hd__a221o_1
X_08283_ net132 net67 net1640 VGND VGND VPWR VPWR _05425_ sky130_fd_sc_hd__mux2_1
Xclkload8 clknet_5_17__leaf_clk VGND VGND VPWR VPWR clkload8/Y sky130_fd_sc_hd__inv_6
XFILLER_165_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07234_ data_array.data0\[1\]\[45\] net1535 net1439 data_array.data0\[2\]\[45\] VGND
+ VGND VPWR VPWR _04494_ sky130_fd_sc_hd__a22o_1
X_07165_ _04430_ _04431_ VGND VGND VPWR VPWR _00031_ sky130_fd_sc_hd__or2_1
XFILLER_118_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06116_ data_array.rdata0\[31\] net1140 net1114 data_array.rdata1\[31\] VGND VGND
+ VPWR VPWR net287 sky130_fd_sc_hd__a22o_1
XFILLER_161_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07096_ data_array.data0\[4\]\[32\] net1330 net1236 data_array.data0\[7\]\[32\] _04368_
+ VGND VGND VPWR VPWR _04369_ sky130_fd_sc_hd__a221o_1
XFILLER_160_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06047_ net1158 net5 fsm.tag_out1\[6\] net1131 VGND VGND VPWR VPWR _03487_ sky130_fd_sc_hd__a22o_1
XFILLER_182_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_184_3886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_184_3897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09806_ net987 net2405 net390 VGND VGND VPWR VPWR _01557_ sky130_fd_sc_hd__mux2_1
XFILLER_59_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07998_ data_array.data1\[0\]\[50\] net1337 net1243 data_array.data1\[3\]\[50\] _05188_
+ VGND VGND VPWR VPWR _05189_ sky130_fd_sc_hd__a221o_1
XFILLER_46_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09737_ net740 net4419 net684 VGND VGND VPWR VPWR _01489_ sky130_fd_sc_hd__mux2_1
X_06949_ data_array.data0\[4\]\[19\] net1390 net1296 data_array.data0\[7\]\[19\] _04234_
+ VGND VGND VPWR VPWR _04235_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_2_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_66_clk clknet_5_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_66_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_83_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09668_ net716 net3257 net613 VGND VGND VPWR VPWR _01420_ sky130_fd_sc_hd__mux2_1
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08619_ net746 net2686 net522 VGND VGND VPWR VPWR _00378_ sky130_fd_sc_hd__mux2_1
X_09599_ net955 net4525 net397 VGND VGND VPWR VPWR _01351_ sky130_fd_sc_hd__mux2_1
X_11630_ clknet_leaf_101_clk _00438_ VGND VGND VPWR VPWR tag_array.tag1\[3\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_46_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_554 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11561_ clknet_leaf_31_clk _00369_ VGND VGND VPWR VPWR tag_array.tag1\[5\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_13300_ clknet_leaf_61_clk _01930_ VGND VGND VPWR VPWR data_array.data0\[10\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_10512_ net897 net3519 net344 VGND VGND VPWR VPWR _02257_ sky130_fd_sc_hd__mux2_1
X_14280_ clknet_leaf_174_clk _02909_ VGND VGND VPWR VPWR data_array.data1\[11\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_11492_ clknet_leaf_153_clk _00301_ VGND VGND VPWR VPWR tag_array.valid0\[3\] sky130_fd_sc_hd__dfxtp_1
X_13231_ clknet_leaf_73_clk _01861_ VGND VGND VPWR VPWR data_array.data0\[11\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_10443_ net1858 net883 net662 VGND VGND VPWR VPWR _02189_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_21_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13162_ clknet_leaf_188_clk _01856_ VGND VGND VPWR VPWR tag_array.tag1\[8\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_10374_ net704 net3442 net540 VGND VGND VPWR VPWR _02121_ sky130_fd_sc_hd__mux2_1
XFILLER_108_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12113_ clknet_leaf_41_clk _00921_ VGND VGND VPWR VPWR data_array.data1\[14\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
X_13093_ clknet_leaf_79_clk _01787_ VGND VGND VPWR VPWR data_array.data1\[13\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
X_12044_ clknet_leaf_221_clk _00852_ VGND VGND VPWR VPWR data_array.data0\[6\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_172_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout790 _05367_ VGND VGND VPWR VPWR net790 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13995_ clknet_leaf_255_clk _02624_ VGND VGND VPWR VPWR data_array.data1\[5\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_57_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_57_clk sky130_fd_sc_hd__clkbuf_8
X_12946_ clknet_leaf_25_clk _01640_ VGND VGND VPWR VPWR data_array.data0\[13\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_142_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_66_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12877_ clknet_leaf_27_clk _01571_ VGND VGND VPWR VPWR data_array.data0\[12\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_103_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11828_ clknet_leaf_71_clk _00636_ VGND VGND VPWR VPWR data_array.data0\[7\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_83_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11759_ clknet_leaf_4_clk _00567_ VGND VGND VPWR VPWR data_array.data0\[8\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_159_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14478_ clknet_leaf_124_clk _03101_ VGND VGND VPWR VPWR data_array.data1\[7\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload103 clknet_leaf_38_clk VGND VGND VPWR VPWR clkload103/Y sky130_fd_sc_hd__clkinv_4
Xclkload114 clknet_leaf_97_clk VGND VGND VPWR VPWR clkload114/Y sky130_fd_sc_hd__bufinv_16
Xclkload125 clknet_leaf_80_clk VGND VGND VPWR VPWR clkload125/Y sky130_fd_sc_hd__inv_8
X_13429_ clknet_leaf_56_clk _02059_ VGND VGND VPWR VPWR data_array.data1\[8\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload136 clknet_leaf_218_clk VGND VGND VPWR VPWR clkload136/Y sky130_fd_sc_hd__inv_8
Xclkload147 clknet_leaf_212_clk VGND VGND VPWR VPWR clkload147/Y sky130_fd_sc_hd__clkinv_2
Xclkload158 clknet_leaf_171_clk VGND VGND VPWR VPWR clkload158/X sky130_fd_sc_hd__clkbuf_4
XFILLER_6_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload169 clknet_leaf_193_clk VGND VGND VPWR VPWR clkload169/Y sky130_fd_sc_hd__clkinv_2
XFILLER_142_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08970_ net884 net2835 net427 VGND VGND VPWR VPWR _00726_ sky130_fd_sc_hd__mux2_1
XFILLER_143_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_166_3550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2606 tag_array.tag0\[5\]\[6\] VGND VGND VPWR VPWR net4257 sky130_fd_sc_hd__dlygate4sd3_1
X_07921_ data_array.data1\[4\]\[43\] net1378 net1284 data_array.data1\[7\]\[43\] _05118_
+ VGND VGND VPWR VPWR _05119_ sky130_fd_sc_hd__a221o_1
Xhold2617 tag_array.tag1\[13\]\[14\] VGND VGND VPWR VPWR net4268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2628 data_array.data0\[6\]\[19\] VGND VGND VPWR VPWR net4279 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2639 data_array.data1\[3\]\[50\] VGND VGND VPWR VPWR net4290 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1905 data_array.data1\[7\]\[58\] VGND VGND VPWR VPWR net3556 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_127_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07852_ data_array.data1\[13\]\[37\] net1544 net1448 data_array.data1\[14\]\[37\]
+ VGND VGND VPWR VPWR _05056_ sky130_fd_sc_hd__a22o_1
Xhold1916 data_array.data1\[9\]\[6\] VGND VGND VPWR VPWR net3567 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1927 data_array.data1\[12\]\[62\] VGND VGND VPWR VPWR net3578 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1938 data_array.data0\[8\]\[39\] VGND VGND VPWR VPWR net3589 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_162_3469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06803_ data_array.data0\[9\]\[6\] net1522 net1426 data_array.data0\[10\]\[6\] VGND
+ VGND VPWR VPWR _04102_ sky130_fd_sc_hd__a22o_1
Xhold1949 data_array.data0\[15\]\[43\] VGND VGND VPWR VPWR net3600 sky130_fd_sc_hd__dlygate4sd3_1
Xinput1 cpu_addr[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
X_07783_ data_array.data1\[12\]\[31\] net1384 net1290 data_array.data1\[15\]\[31\]
+ _04992_ VGND VGND VPWR VPWR _04993_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_48_clk clknet_5_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_48_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_37_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09522_ net739 net3326 net623 VGND VGND VPWR VPWR _01275_ sky130_fd_sc_hd__mux2_1
X_06734_ net1196 _04033_ _04037_ net1622 VGND VGND VPWR VPWR _04040_ sky130_fd_sc_hd__a22o_1
XFILLER_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09453_ net820 net3457 _05570_ VGND VGND VPWR VPWR _01206_ sky130_fd_sc_hd__mux2_1
XFILLER_149_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06665_ tag_array.tag1\[8\]\[18\] net1372 net1278 tag_array.tag1\[11\]\[18\] _03976_
+ VGND VGND VPWR VPWR _03977_ sky130_fd_sc_hd__a221o_1
XFILLER_169_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08404_ net1128 _05505_ VGND VGND VPWR VPWR _05506_ sky130_fd_sc_hd__and2_1
X_05616_ fsm.tag_out1\[6\] VGND VGND VPWR VPWR _03138_ sky130_fd_sc_hd__inv_2
X_09384_ net866 net2810 net405 VGND VGND VPWR VPWR _01137_ sky130_fd_sc_hd__mux2_1
X_06596_ tag_array.tag1\[5\]\[12\] net1592 net1496 tag_array.tag1\[6\]\[12\] VGND
+ VGND VPWR VPWR _03914_ sky130_fd_sc_hd__a22o_1
X_08335_ net1129 _05459_ VGND VGND VPWR VPWR _05460_ sky130_fd_sc_hd__and2_1
XFILLER_177_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08266_ net163 net1159 net25 VGND VGND VPWR VPWR _05412_ sky130_fd_sc_hd__and3_1
XFILLER_20_596 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07217_ data_array.data0\[4\]\[43\] net1377 net1283 data_array.data0\[7\]\[43\] _04478_
+ VGND VGND VPWR VPWR _04479_ sky130_fd_sc_hd__a221o_1
XFILLER_153_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08197_ _03135_ _03147_ VGND VGND VPWR VPWR _05366_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_18_Left_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_996 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07148_ data_array.data0\[13\]\[37\] net1547 net1451 data_array.data0\[14\]\[37\]
+ VGND VGND VPWR VPWR _04416_ sky130_fd_sc_hd__a22o_1
XFILLER_180_549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07079_ data_array.data0\[12\]\[31\] net1385 net1291 data_array.data0\[15\]\[31\]
+ _04352_ VGND VGND VPWR VPWR _04353_ sky130_fd_sc_hd__a221o_1
XFILLER_161_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_55 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10090_ net3505 net765 net642 VGND VGND VPWR VPWR _01839_ sky130_fd_sc_hd__mux2_1
Xfanout1007 _05472_ VGND VGND VPWR VPWR net1007 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_160_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1018 _05466_ VGND VGND VPWR VPWR net1018 sky130_fd_sc_hd__clkbuf_2
Xfanout1029 _05460_ VGND VGND VPWR VPWR net1029 sky130_fd_sc_hd__buf_1
XFILLER_99_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_27_Left_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_39_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_39_clk sky130_fd_sc_hd__clkbuf_8
X_12800_ clknet_leaf_186_clk _01494_ VGND VGND VPWR VPWR tag_array.tag1\[10\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_48_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13780_ clknet_leaf_85_clk _02409_ VGND VGND VPWR VPWR data_array.data1\[2\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_10992_ net1734 net1032 net341 VGND VGND VPWR VPWR _02736_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12731_ clknet_leaf_190_clk _01425_ VGND VGND VPWR VPWR tag_array.tag0\[7\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12662_ clknet_leaf_84_clk _01356_ VGND VGND VPWR VPWR data_array.data0\[15\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14401_ clknet_leaf_5_clk _03024_ VGND VGND VPWR VPWR data_array.data1\[10\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
X_11613_ clknet_leaf_194_clk _00421_ VGND VGND VPWR VPWR tag_array.tag1\[3\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12593_ clknet_leaf_106_clk _01287_ VGND VGND VPWR VPWR tag_array.tag0\[0\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_169_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14332_ clknet_leaf_212_clk _02961_ VGND VGND VPWR VPWR data_array.data1\[11\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
X_11544_ clknet_leaf_103_clk _00352_ VGND VGND VPWR VPWR tag_array.tag1\[6\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_36_Left_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14263_ clknet_leaf_77_clk _02892_ VGND VGND VPWR VPWR data_array.data1\[12\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_1041 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11475_ clknet_leaf_172_clk _00285_ VGND VGND VPWR VPWR tag_array.valid1\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_143_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13214_ clknet_leaf_2_clk _00110_ VGND VGND VPWR VPWR data_array.rdata1\[51\] sky130_fd_sc_hd__dfxtp_1
X_10426_ net2735 net950 net671 VGND VGND VPWR VPWR _02172_ sky130_fd_sc_hd__mux2_1
X_14194_ clknet_leaf_93_clk _02823_ VGND VGND VPWR VPWR data_array.data0\[2\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_100_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13145_ clknet_leaf_134_clk _01839_ VGND VGND VPWR VPWR tag_array.tag1\[8\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_125_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10357_ net770 net2887 net540 VGND VGND VPWR VPWR _02104_ sky130_fd_sc_hd__mux2_1
X_13076_ clknet_leaf_248_clk _01770_ VGND VGND VPWR VPWR data_array.data1\[13\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_10288_ net2021 net1011 net633 VGND VGND VPWR VPWR _02035_ sky130_fd_sc_hd__mux2_1
XFILLER_105_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12027_ clknet_leaf_216_clk _00835_ VGND VGND VPWR VPWR data_array.data0\[6\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout1530 net1543 VGND VGND VPWR VPWR net1530 sky130_fd_sc_hd__clkbuf_2
XFILLER_111_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1541 net1542 VGND VGND VPWR VPWR net1541 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_144_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1552 net1554 VGND VGND VPWR VPWR net1552 sky130_fd_sc_hd__clkbuf_4
Xfanout1563 net1566 VGND VGND VPWR VPWR net1563 sky130_fd_sc_hd__clkbuf_2
XFILLER_66_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_45_Left_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1574 net1576 VGND VGND VPWR VPWR net1574 sky130_fd_sc_hd__clkbuf_4
Xfanout1585 net1587 VGND VGND VPWR VPWR net1585 sky130_fd_sc_hd__clkbuf_4
Xfanout1596 net1613 VGND VGND VPWR VPWR net1596 sky130_fd_sc_hd__clkbuf_4
XFILLER_53_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13978_ clknet_leaf_18_clk _02607_ VGND VGND VPWR VPWR data_array.data1\[5\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12929_ clknet_leaf_72_clk _01623_ VGND VGND VPWR VPWR data_array.data0\[13\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_73_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06450_ _03780_ _03781_ VGND VGND VPWR VPWR _00146_ sky130_fd_sc_hd__or2_1
X_06381_ tag_array.tag0\[0\]\[17\] net1412 net1318 tag_array.tag0\[3\]\[17\] _03718_
+ VGND VGND VPWR VPWR _03719_ sky130_fd_sc_hd__a221o_1
XFILLER_147_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08120_ net1196 _05293_ _05297_ net1622 VGND VGND VPWR VPWR _05300_ sky130_fd_sc_hd__a22o_1
XFILLER_119_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08051_ data_array.data1\[8\]\[55\] net1344 net1250 data_array.data1\[11\]\[55\]
+ _05236_ VGND VGND VPWR VPWR _05237_ sky130_fd_sc_hd__a221o_1
XFILLER_119_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07002_ data_array.data0\[12\]\[24\] net1385 net1291 data_array.data0\[15\]\[24\]
+ _04282_ VGND VGND VPWR VPWR _04283_ sky130_fd_sc_hd__a221o_1
XFILLER_179_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_164_3509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08953_ net954 net2769 net429 VGND VGND VPWR VPWR _00709_ sky130_fd_sc_hd__mux2_1
Xhold2403 data_array.data1\[5\]\[11\] VGND VGND VPWR VPWR net4054 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2414 data_array.data0\[14\]\[44\] VGND VGND VPWR VPWR net4065 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_181_3834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2425 tag_array.tag0\[11\]\[15\] VGND VGND VPWR VPWR net4076 sky130_fd_sc_hd__dlygate4sd3_1
X_07904_ data_array.data1\[8\]\[42\] net1396 net1302 data_array.data1\[11\]\[42\]
+ _05102_ VGND VGND VPWR VPWR _05103_ sky130_fd_sc_hd__a221o_1
Xhold2436 data_array.data0\[12\]\[54\] VGND VGND VPWR VPWR net4087 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_181_3845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1702 data_array.data0\[5\]\[0\] VGND VGND VPWR VPWR net3353 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_1051 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08884_ net971 net4162 net434 VGND VGND VPWR VPWR _00641_ sky130_fd_sc_hd__mux2_1
Xhold2447 data_array.data1\[3\]\[12\] VGND VGND VPWR VPWR net4098 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2458 data_array.data1\[9\]\[23\] VGND VGND VPWR VPWR net4109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1713 tag_array.tag1\[4\]\[3\] VGND VGND VPWR VPWR net3364 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1724 data_array.data0\[9\]\[38\] VGND VGND VPWR VPWR net3375 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2469 tag_array.tag0\[13\]\[4\] VGND VGND VPWR VPWR net4120 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1735 tag_array.tag1\[7\]\[14\] VGND VGND VPWR VPWR net3386 sky130_fd_sc_hd__dlygate4sd3_1
X_07835_ net1166 _05035_ _05039_ net1214 VGND VGND VPWR VPWR _05041_ sky130_fd_sc_hd__a22o_1
XFILLER_84_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1746 data_array.data0\[1\]\[7\] VGND VGND VPWR VPWR net3397 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1757 data_array.data0\[13\]\[42\] VGND VGND VPWR VPWR net3408 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1768 data_array.data0\[15\]\[34\] VGND VGND VPWR VPWR net3419 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1779 tag_array.tag0\[2\]\[9\] VGND VGND VPWR VPWR net3430 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07766_ data_array.data1\[5\]\[29\] net1572 net1476 data_array.data1\[6\]\[29\] VGND
+ VGND VPWR VPWR _04978_ sky130_fd_sc_hd__a22o_1
XFILLER_84_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09505_ net709 net3229 net625 VGND VGND VPWR VPWR _01258_ sky130_fd_sc_hd__mux2_1
XFILLER_112_46 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06717_ tag_array.tag1\[5\]\[23\] net1610 net1514 tag_array.tag1\[6\]\[23\] VGND
+ VGND VPWR VPWR _04024_ sky130_fd_sc_hd__a22o_1
X_07697_ data_array.data1\[0\]\[23\] net1359 net1265 data_array.data1\[3\]\[23\] _04914_
+ VGND VGND VPWR VPWR _04915_ sky130_fd_sc_hd__a221o_1
XFILLER_80_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_179_3796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09436_ net923 net2664 net587 VGND VGND VPWR VPWR _01189_ sky130_fd_sc_hd__mux2_1
X_06648_ _03960_ _03961_ VGND VGND VPWR VPWR _00163_ sky130_fd_sc_hd__or2_1
XFILLER_12_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09367_ net933 net4065 net408 VGND VGND VPWR VPWR _01120_ sky130_fd_sc_hd__mux2_1
X_06579_ tag_array.tag1\[4\]\[10\] net1404 net1310 tag_array.tag1\[7\]\[10\] _03898_
+ VGND VGND VPWR VPWR _03899_ sky130_fd_sc_hd__a221o_1
XFILLER_123_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08318_ net1997 net1052 net692 VGND VGND VPWR VPWR _00235_ sky130_fd_sc_hd__mux2_1
XFILLER_162_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_50 net806 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09298_ net788 net3343 net544 VGND VGND VPWR VPWR _01052_ sky130_fd_sc_hd__mux2_1
XFILLER_165_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_61 net1495 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_72 _03127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_83 net1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08249_ fsm.tag_out1\[18\] net816 net808 fsm.tag_out0\[18\] _05400_ VGND VGND VPWR
+ VPWR _05401_ sky130_fd_sc_hd__a221o_1
XFILLER_153_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11260_ net991 net4411 net681 VGND VGND VPWR VPWR _03003_ sky130_fd_sc_hd__mux2_1
XFILLER_180_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10211_ net962 net2802 net357 VGND VGND VPWR VPWR _01958_ sky130_fd_sc_hd__mux2_1
XFILLER_133_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11191_ net1011 net4299 net648 VGND VGND VPWR VPWR _02934_ sky130_fd_sc_hd__mux2_1
XFILLER_107_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10142_ net976 net3921 net367 VGND VGND VPWR VPWR _01890_ sky130_fd_sc_hd__mux2_1
Xoutput190 net190 VGND VGND VPWR VPWR cpu_rdata[32] sky130_fd_sc_hd__buf_4
X_10073_ net732 net3212 net599 VGND VGND VPWR VPWR _01822_ sky130_fd_sc_hd__mux2_1
XFILLER_75_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2970 data_array.data0\[10\]\[1\] VGND VGND VPWR VPWR net4621 sky130_fd_sc_hd__dlygate4sd3_1
X_13901_ clknet_leaf_198_clk _02530_ VGND VGND VPWR VPWR data_array.data1\[4\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_153_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13832_ clknet_leaf_174_clk _02461_ VGND VGND VPWR VPWR data_array.data1\[3\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13763_ clknet_leaf_55_clk _02392_ VGND VGND VPWR VPWR data_array.data1\[1\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
X_10975_ net2550 net1102 net339 VGND VGND VPWR VPWR _02719_ sky130_fd_sc_hd__mux2_1
XFILLER_55_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12714_ clknet_leaf_143_clk _01408_ VGND VGND VPWR VPWR tag_array.tag0\[7\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_13694_ clknet_leaf_216_clk _02323_ VGND VGND VPWR VPWR data_array.data1\[15\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_80_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_0__f_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_5_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_80_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12645_ clknet_leaf_237_clk _01339_ VGND VGND VPWR VPWR data_array.data0\[15\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12576_ clknet_leaf_137_clk _01270_ VGND VGND VPWR VPWR tag_array.tag0\[10\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_178_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_866 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14315_ clknet_leaf_259_clk _02944_ VGND VGND VPWR VPWR data_array.data1\[11\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11527_ clknet_leaf_174_clk _00335_ VGND VGND VPWR VPWR tag_array.valid1\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_156_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14246_ clknet_leaf_68_clk _02875_ VGND VGND VPWR VPWR data_array.data1\[12\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold309 data_array.data1\[4\]\[42\] VGND VGND VPWR VPWR net1960 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11458_ clknet_leaf_91_clk _00268_ VGND VGND VPWR VPWR data_array.data0\[0\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_172_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10409_ net2149 net1016 net664 VGND VGND VPWR VPWR _02155_ sky130_fd_sc_hd__mux2_1
X_14177_ clknet_leaf_0_clk _02806_ VGND VGND VPWR VPWR data_array.data0\[2\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_11389_ clknet_leaf_191_clk _00199_ VGND VGND VPWR VPWR tag_array.tag1\[7\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_112_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13128_ clknet_leaf_164_clk _01822_ VGND VGND VPWR VPWR tag_array.tag0\[3\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_13059_ clknet_leaf_119_clk _01753_ VGND VGND VPWR VPWR data_array.data1\[13\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_05950_ net131 net1151 _03426_ _03427_ VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__a22o_1
XFILLER_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1009 data_array.data1\[5\]\[8\] VGND VGND VPWR VPWR net2660 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1360 net1364 VGND VGND VPWR VPWR net1360 sky130_fd_sc_hd__clkbuf_4
XFILLER_38_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1371 net1375 VGND VGND VPWR VPWR net1371 sky130_fd_sc_hd__clkbuf_4
X_05881_ net106 net1152 _03380_ _03381_ VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__a22o_1
XFILLER_38_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1382 net1383 VGND VGND VPWR VPWR net1382 sky130_fd_sc_hd__clkbuf_2
Xfanout1393 net1394 VGND VGND VPWR VPWR net1393 sky130_fd_sc_hd__clkbuf_4
X_07620_ data_array.data1\[4\]\[16\] net1354 net1260 data_array.data1\[7\]\[16\] _04844_
+ VGND VGND VPWR VPWR _04845_ sky130_fd_sc_hd__a221o_1
XFILLER_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_886 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07551_ data_array.data1\[9\]\[10\] net1606 net1510 data_array.data1\[10\]\[10\]
+ VGND VGND VPWR VPWR _04782_ sky130_fd_sc_hd__a22o_1
XFILLER_35_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06502_ tag_array.tag1\[0\]\[3\] net1361 net1267 tag_array.tag1\[3\]\[3\] _03828_
+ VGND VGND VPWR VPWR _03829_ sky130_fd_sc_hd__a221o_1
X_07482_ net1194 _04713_ _04717_ net1620 VGND VGND VPWR VPWR _04720_ sky130_fd_sc_hd__a22o_1
X_09221_ net696 net2805 net632 VGND VGND VPWR VPWR _00975_ sky130_fd_sc_hd__mux2_1
X_06433_ tag_array.tag0\[13\]\[22\] net1565 net1469 tag_array.tag0\[14\]\[22\] VGND
+ VGND VPWR VPWR _03766_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_157_3379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09152_ net935 net3198 net575 VGND VGND VPWR VPWR _00906_ sky130_fd_sc_hd__mux2_1
X_06364_ tag_array.tag0\[8\]\[16\] net1409 net1315 tag_array.tag0\[11\]\[16\] _03702_
+ VGND VGND VPWR VPWR _03703_ sky130_fd_sc_hd__a221o_1
X_08103_ data_array.data1\[5\]\[60\] net1604 net1508 data_array.data1\[6\]\[60\] VGND
+ VGND VPWR VPWR _05284_ sky130_fd_sc_hd__a22o_1
X_09083_ net954 net2324 net413 VGND VGND VPWR VPWR _00837_ sky130_fd_sc_hd__mux2_1
X_06295_ net1230 _03635_ _03639_ net1182 VGND VGND VPWR VPWR _03641_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_135_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08034_ _05220_ _05221_ VGND VGND VPWR VPWR _00112_ sky130_fd_sc_hd__or2_1
Xinput70 cpu_wdata[42] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_1
Xhold810 data_array.data0\[7\]\[17\] VGND VGND VPWR VPWR net2461 sky130_fd_sc_hd__dlygate4sd3_1
Xinput81 cpu_wdata[52] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_1
Xhold821 data_array.data0\[2\]\[33\] VGND VGND VPWR VPWR net2472 sky130_fd_sc_hd__dlygate4sd3_1
Xinput92 cpu_wdata[62] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_1
Xhold832 data_array.data1\[9\]\[8\] VGND VGND VPWR VPWR net2483 sky130_fd_sc_hd__dlygate4sd3_1
Xhold843 data_array.data1\[9\]\[27\] VGND VGND VPWR VPWR net2494 sky130_fd_sc_hd__dlygate4sd3_1
Xhold854 data_array.data0\[2\]\[4\] VGND VGND VPWR VPWR net2505 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold865 tag_array.tag1\[12\]\[0\] VGND VGND VPWR VPWR net2516 sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 data_array.data0\[2\]\[34\] VGND VGND VPWR VPWR net2527 sky130_fd_sc_hd__dlygate4sd3_1
Xhold887 data_array.data0\[4\]\[57\] VGND VGND VPWR VPWR net2538 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_107_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold898 data_array.data1\[10\]\[15\] VGND VGND VPWR VPWR net2549 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_107_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09985_ net888 net4437 net371 VGND VGND VPWR VPWR _01734_ sky130_fd_sc_hd__mux2_1
XFILLER_89_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2200 data_array.data0\[6\]\[48\] VGND VGND VPWR VPWR net3851 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2211 data_array.data1\[7\]\[34\] VGND VGND VPWR VPWR net3862 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2222 data_array.data1\[6\]\[35\] VGND VGND VPWR VPWR net3873 sky130_fd_sc_hd__dlygate4sd3_1
X_08936_ net1020 net2906 net427 VGND VGND VPWR VPWR _00692_ sky130_fd_sc_hd__mux2_1
Xhold2233 data_array.data0\[14\]\[0\] VGND VGND VPWR VPWR net3884 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_36_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2244 data_array.data1\[5\]\[9\] VGND VGND VPWR VPWR net3895 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2255 data_array.data1\[7\]\[42\] VGND VGND VPWR VPWR net3906 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1510 data_array.data0\[13\]\[31\] VGND VGND VPWR VPWR net3161 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1521 data_array.data0\[13\]\[39\] VGND VGND VPWR VPWR net3172 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2266 data_array.data1\[12\]\[50\] VGND VGND VPWR VPWR net3917 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08867_ net1036 net4226 net439 VGND VGND VPWR VPWR _00624_ sky130_fd_sc_hd__mux2_1
Xhold1532 tag_array.tag1\[3\]\[11\] VGND VGND VPWR VPWR net3183 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2277 data_array.data1\[1\]\[29\] VGND VGND VPWR VPWR net3928 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2288 tag_array.tag1\[10\]\[6\] VGND VGND VPWR VPWR net3939 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1543 data_array.data0\[9\]\[47\] VGND VGND VPWR VPWR net3194 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2299 data_array.data0\[14\]\[48\] VGND VGND VPWR VPWR net3950 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1554 data_array.data0\[15\]\[7\] VGND VGND VPWR VPWR net3205 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1565 tag_array.tag1\[9\]\[10\] VGND VGND VPWR VPWR net3216 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1576 data_array.data0\[8\]\[1\] VGND VGND VPWR VPWR net3227 sky130_fd_sc_hd__dlygate4sd3_1
X_07818_ data_array.data1\[4\]\[34\] net1340 net1246 data_array.data1\[7\]\[34\] _05024_
+ VGND VGND VPWR VPWR _05025_ sky130_fd_sc_hd__a221o_1
XFILLER_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1587 data_array.data0\[7\]\[15\] VGND VGND VPWR VPWR net3238 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_28_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08798_ net2006 net1052 net446 VGND VGND VPWR VPWR _00556_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1598 data_array.data1\[9\]\[43\] VGND VGND VPWR VPWR net3249 sky130_fd_sc_hd__dlygate4sd3_1
X_07749_ data_array.data1\[9\]\[28\] net1541 net1445 data_array.data1\[10\]\[28\]
+ VGND VGND VPWR VPWR _04962_ sky130_fd_sc_hd__a22o_1
X_10760_ net934 net3775 net498 VGND VGND VPWR VPWR _02505_ sky130_fd_sc_hd__mux2_1
XFILLER_16_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09419_ net990 net3300 net586 VGND VGND VPWR VPWR _01172_ sky130_fd_sc_hd__mux2_1
X_10691_ net1947 net952 net479 VGND VGND VPWR VPWR _02436_ sky130_fd_sc_hd__mux2_1
XFILLER_12_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12430_ clknet_leaf_57_clk _01124_ VGND VGND VPWR VPWR data_array.data0\[14\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12361_ clknet_leaf_49_clk _00037_ VGND VGND VPWR VPWR data_array.rdata0\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14100_ clknet_leaf_94_clk _02729_ VGND VGND VPWR VPWR data_array.data0\[1\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_11312_ net1044 net3390 net798 VGND VGND VPWR VPWR _03055_ sky130_fd_sc_hd__mux2_1
XFILLER_126_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12292_ clknet_leaf_188_clk _01050_ VGND VGND VPWR VPWR tag_array.tag1\[13\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14031_ clknet_leaf_82_clk _02660_ VGND VGND VPWR VPWR data_array.data1\[6\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_11243_ net1057 net2112 net677 VGND VGND VPWR VPWR _02986_ sky130_fd_sc_hd__mux2_1
XFILLER_164_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11174_ net1079 net2918 net650 VGND VGND VPWR VPWR _02917_ sky130_fd_sc_hd__mux2_1
XFILLER_161_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_270_clk clknet_5_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_270_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10125_ net1046 net3331 net364 VGND VGND VPWR VPWR _01873_ sky130_fd_sc_hd__mux2_1
XFILLER_67_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10056_ net863 net2559 net564 VGND VGND VPWR VPWR _01805_ sky130_fd_sc_hd__mux2_1
XFILLER_57_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13815_ clknet_leaf_78_clk _02444_ VGND VGND VPWR VPWR data_array.data1\[2\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_169_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13746_ clknet_leaf_88_clk _02375_ VGND VGND VPWR VPWR data_array.data1\[1\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
X_10958_ net908 net3723 net526 VGND VGND VPWR VPWR _02703_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_139_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13677_ clknet_leaf_217_clk _02306_ VGND VGND VPWR VPWR data_array.data1\[15\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_176_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10889_ net930 net3414 net518 VGND VGND VPWR VPWR _02634_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12628_ clknet_leaf_111_clk _01322_ VGND VGND VPWR VPWR data_array.data0\[15\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_117_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12559_ clknet_leaf_157_clk _01253_ VGND VGND VPWR VPWR tag_array.tag0\[11\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_157_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06080_ fsm.tag_out0\[22\] net1120 _03503_ VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__a21o_1
Xhold106 data_array.data1\[8\]\[26\] VGND VGND VPWR VPWR net1757 sky130_fd_sc_hd__dlygate4sd3_1
Xhold117 data_array.data0\[8\]\[45\] VGND VGND VPWR VPWR net1768 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold128 data_array.data1\[4\]\[45\] VGND VGND VPWR VPWR net1779 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold139 data_array.data1\[4\]\[47\] VGND VGND VPWR VPWR net1790 sky130_fd_sc_hd__dlygate4sd3_1
X_14229_ clknet_leaf_199_clk _02858_ VGND VGND VPWR VPWR data_array.data1\[12\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_508 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_130_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout608 _05579_ VGND VGND VPWR VPWR net608 sky130_fd_sc_hd__buf_2
XFILLER_112_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout619 net620 VGND VGND VPWR VPWR net619 sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_261_clk clknet_5_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_261_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_98_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_107_Right_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09770_ net1934 net706 net672 VGND VGND VPWR VPWR _01522_ sky130_fd_sc_hd__mux2_1
X_06982_ data_array.data0\[0\]\[22\] net1341 net1247 data_array.data0\[3\]\[22\] _04264_
+ VGND VGND VPWR VPWR _04265_ sky130_fd_sc_hd__a221o_1
XFILLER_86_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08721_ net2142 net740 net476 VGND VGND VPWR VPWR _00480_ sky130_fd_sc_hd__mux2_1
X_05933_ data_array.rdata0\[34\] net847 net1143 VGND VGND VPWR VPWR _03416_ sky130_fd_sc_hd__o21a_1
XFILLER_100_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1190 net1191 VGND VGND VPWR VPWR net1190 sky130_fd_sc_hd__buf_4
XFILLER_67_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08652_ net1817 net714 net512 VGND VGND VPWR VPWR _00411_ sky130_fd_sc_hd__mux2_1
X_05864_ net851 data_array.rdata0\[11\] net1148 VGND VGND VPWR VPWR _03370_ sky130_fd_sc_hd__o21a_1
XFILLER_93_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07603_ net1628 _04823_ _04827_ net1202 VGND VGND VPWR VPWR _04830_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_159_3419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08583_ net791 net3135 net531 VGND VGND VPWR VPWR _00342_ sky130_fd_sc_hd__mux2_1
XFILLER_54_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05795_ fsm.tag_out1\[19\] net19 VGND VGND VPWR VPWR _03312_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_176_3733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07534_ data_array.data1\[8\]\[8\] net1345 net1251 data_array.data1\[11\]\[8\] _04766_
+ VGND VGND VPWR VPWR _04767_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_176_3744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07465_ data_array.data1\[5\]\[2\] net1530 net1434 data_array.data1\[6\]\[2\] VGND
+ VGND VPWR VPWR _04704_ sky130_fd_sc_hd__a22o_1
X_09204_ net762 net2099 net632 VGND VGND VPWR VPWR _00958_ sky130_fd_sc_hd__mux2_1
X_06416_ net1173 _03745_ _03749_ net1222 VGND VGND VPWR VPWR _03751_ sky130_fd_sc_hd__a22o_1
XFILLER_167_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07396_ _04640_ _04641_ VGND VGND VPWR VPWR _00054_ sky130_fd_sc_hd__or2_1
XFILLER_176_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09135_ net1001 net3643 net567 VGND VGND VPWR VPWR _00889_ sky130_fd_sc_hd__mux2_1
X_06347_ tag_array.tag0\[1\]\[14\] net1558 net1462 tag_array.tag0\[2\]\[14\] VGND
+ VGND VPWR VPWR _03688_ sky130_fd_sc_hd__a22o_1
XFILLER_33_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09066_ net1020 net4177 net411 VGND VGND VPWR VPWR _00820_ sky130_fd_sc_hd__mux2_1
XFILLER_108_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06278_ tag_array.tag0\[0\]\[8\] net1410 net1316 tag_array.tag0\[3\]\[8\] _03624_
+ VGND VGND VPWR VPWR _03625_ sky130_fd_sc_hd__a221o_1
X_08017_ data_array.data1\[9\]\[52\] net1545 net1449 data_array.data1\[10\]\[52\]
+ VGND VGND VPWR VPWR _05206_ sky130_fd_sc_hd__a22o_1
XFILLER_151_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold640 data_array.data1\[14\]\[58\] VGND VGND VPWR VPWR net2291 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold651 data_array.data0\[6\]\[62\] VGND VGND VPWR VPWR net2302 sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 data_array.data0\[11\]\[12\] VGND VGND VPWR VPWR net2313 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold673 data_array.data0\[6\]\[39\] VGND VGND VPWR VPWR net2324 sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 data_array.data1\[6\]\[19\] VGND VGND VPWR VPWR net2335 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold695 data_array.data1\[5\]\[43\] VGND VGND VPWR VPWR net2346 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_252_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_252_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_34_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09968_ net956 net4269 net375 VGND VGND VPWR VPWR _01717_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_34_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2030 data_array.data0\[9\]\[22\] VGND VGND VPWR VPWR net3681 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2041 data_array.data1\[9\]\[53\] VGND VGND VPWR VPWR net3692 sky130_fd_sc_hd__dlygate4sd3_1
X_08919_ net1088 net3446 net428 VGND VGND VPWR VPWR _00675_ sky130_fd_sc_hd__mux2_1
Xhold2052 tag_array.tag0\[0\]\[7\] VGND VGND VPWR VPWR net3703 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2063 tag_array.tag0\[7\]\[3\] VGND VGND VPWR VPWR net3714 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09899_ net873 net4396 net382 VGND VGND VPWR VPWR _01649_ sky130_fd_sc_hd__mux2_1
Xhold2074 data_array.data1\[9\]\[24\] VGND VGND VPWR VPWR net3725 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_40_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1340 data_array.data1\[15\]\[21\] VGND VGND VPWR VPWR net2991 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2085 data_array.data1\[9\]\[29\] VGND VGND VPWR VPWR net3736 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1351 data_array.data0\[5\]\[2\] VGND VGND VPWR VPWR net3002 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2096 tag_array.tag0\[3\]\[9\] VGND VGND VPWR VPWR net3747 sky130_fd_sc_hd__dlygate4sd3_1
X_11930_ clknet_leaf_72_clk _00738_ VGND VGND VPWR VPWR data_array.data0\[4\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1362 tag_array.tag1\[12\]\[21\] VGND VGND VPWR VPWR net3013 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_40_1059 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1373 data_array.data0\[6\]\[8\] VGND VGND VPWR VPWR net3024 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_175_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1384 data_array.data0\[13\]\[35\] VGND VGND VPWR VPWR net3035 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1395 tag_array.tag0\[3\]\[0\] VGND VGND VPWR VPWR net3046 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11861_ clknet_leaf_226_clk _00669_ VGND VGND VPWR VPWR data_array.data0\[7\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_45_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13600_ clknet_leaf_4_clk _02229_ VGND VGND VPWR VPWR data_array.data0\[9\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10812_ net1963 net980 net502 VGND VGND VPWR VPWR _02557_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11792_ clknet_leaf_207_clk _00600_ VGND VGND VPWR VPWR data_array.data0\[8\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_25_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13531_ clknet_leaf_234_clk _02160_ VGND VGND VPWR VPWR data_array.data1\[0\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_10743_ net1000 net3769 net491 VGND VGND VPWR VPWR _02488_ sky130_fd_sc_hd__mux2_1
XFILLER_159_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13462_ clknet_leaf_180_clk _02092_ VGND VGND VPWR VPWR tag_array.tag0\[1\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_159_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10674_ net1849 net1022 net479 VGND VGND VPWR VPWR _02419_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12413_ clknet_leaf_38_clk _01107_ VGND VGND VPWR VPWR data_array.data0\[14\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_13393_ clknet_leaf_199_clk _02023_ VGND VGND VPWR VPWR data_array.data1\[8\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_166_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12344_ clknet_leaf_254_clk _00018_ VGND VGND VPWR VPWR data_array.rdata0\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12275_ clknet_leaf_132_clk _01033_ VGND VGND VPWR VPWR tag_array.tag1\[13\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14014_ clknet_leaf_215_clk _02643_ VGND VGND VPWR VPWR data_array.data1\[5\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
X_11226_ net871 net2453 net658 VGND VGND VPWR VPWR _02969_ sky130_fd_sc_hd__mux2_1
XFILLER_136_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_243_clk clknet_5_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_243_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_71_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11157_ net891 net3780 net543 VGND VGND VPWR VPWR _02900_ sky130_fd_sc_hd__mux2_1
XFILLER_150_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10108_ _05414_ _05550_ VGND VGND VPWR VPWR _03128_ sky130_fd_sc_hd__or2_1
X_11088_ net1775 net910 net329 VGND VGND VPWR VPWR _02831_ sky130_fd_sc_hd__mux2_1
X_10039_ net931 net3679 net556 VGND VGND VPWR VPWR _01788_ sky130_fd_sc_hd__mux2_1
XFILLER_76_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13729_ clknet_leaf_267_clk _02358_ VGND VGND VPWR VPWR data_array.data1\[1\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_154_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07250_ data_array.data0\[0\]\[46\] net1341 net1247 data_array.data0\[3\]\[46\] _04508_
+ VGND VGND VPWR VPWR _04509_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_171_3641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_171_3652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06201_ tag_array.tag0\[4\]\[1\] net1402 net1308 tag_array.tag0\[7\]\[1\] _03554_
+ VGND VGND VPWR VPWR _03555_ sky130_fd_sc_hd__a221o_1
XFILLER_164_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07181_ data_array.data0\[9\]\[40\] net1605 net1509 data_array.data0\[10\]\[40\]
+ VGND VGND VPWR VPWR _04446_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_30_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06132_ data_array.rdata0\[47\] net1139 net1115 data_array.rdata1\[47\] VGND VGND
+ VPWR VPWR net304 sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_132_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06063_ net1158 net14 fsm.tag_out1\[14\] net1131 VGND VGND VPWR VPWR _03495_ sky130_fd_sc_hd__a22o_1
Xfanout405 net409 VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__buf_4
XFILLER_113_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout416 net417 VGND VGND VPWR VPWR net416 sky130_fd_sc_hd__buf_4
XFILLER_59_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout427 net433 VGND VGND VPWR VPWR net427 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_234_clk clknet_5_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_234_clk
+ sky130_fd_sc_hd__clkbuf_8
X_09822_ net920 net2850 net390 VGND VGND VPWR VPWR _01573_ sky130_fd_sc_hd__mux2_1
Xfanout438 net439 VGND VGND VPWR VPWR net438 sky130_fd_sc_hd__buf_4
Xfanout449 _05607_ VGND VGND VPWR VPWR net449 sky130_fd_sc_hd__clkbuf_8
XFILLER_58_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09753_ net2248 net774 net664 VGND VGND VPWR VPWR _01505_ sky130_fd_sc_hd__mux2_1
X_06965_ net1210 _04243_ _04247_ net1636 VGND VGND VPWR VPWR _04250_ sky130_fd_sc_hd__a22o_1
X_08704_ net2103 net706 net488 VGND VGND VPWR VPWR _00463_ sky130_fd_sc_hd__mux2_1
X_05916_ data_array.rdata1\[28\] net829 net838 VGND VGND VPWR VPWR _03405_ sky130_fd_sc_hd__a21o_1
XFILLER_55_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09684_ net752 net2695 net606 VGND VGND VPWR VPWR _01436_ sky130_fd_sc_hd__mux2_1
X_06896_ data_array.data0\[12\]\[14\] net1379 net1285 data_array.data0\[15\]\[14\]
+ _04186_ VGND VGND VPWR VPWR _04187_ sky130_fd_sc_hd__a221o_1
XFILLER_27_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08635_ net1940 net782 net504 VGND VGND VPWR VPWR _00394_ sky130_fd_sc_hd__mux2_1
X_05847_ data_array.rdata1\[5\] net831 net840 VGND VGND VPWR VPWR _03359_ sky130_fd_sc_hd__a21o_1
XFILLER_15_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08566_ net811 _05574_ VGND VGND VPWR VPWR _05598_ sky130_fd_sc_hd__nand2_2
XFILLER_42_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05778_ _03259_ _03264_ _03274_ VGND VGND VPWR VPWR _03295_ sky130_fd_sc_hd__or3_1
X_07517_ _04750_ _04751_ VGND VGND VPWR VPWR _00124_ sky130_fd_sc_hd__or2_1
X_08497_ _03514_ _03519_ net823 VGND VGND VPWR VPWR _05568_ sky130_fd_sc_hd__or3_1
XFILLER_167_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07448_ data_array.data1\[4\]\[0\] net1367 net1272 data_array.data1\[7\]\[0\] _04688_
+ VGND VGND VPWR VPWR _04689_ sky130_fd_sc_hd__a221o_1
XFILLER_11_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07379_ data_array.data0\[13\]\[58\] net1548 net1452 data_array.data0\[14\]\[58\]
+ VGND VGND VPWR VPWR _04626_ sky130_fd_sc_hd__a22o_1
X_09118_ net1070 net2460 net576 VGND VGND VPWR VPWR _00872_ sky130_fd_sc_hd__mux2_1
XFILLER_109_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10390_ net1823 net1094 net668 VGND VGND VPWR VPWR _02136_ sky130_fd_sc_hd__mux2_1
XFILLER_159_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09049_ net1088 net2687 net412 VGND VGND VPWR VPWR _00803_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_92_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_880 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12060_ clknet_leaf_268_clk _00868_ VGND VGND VPWR VPWR data_array.data1\[14\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold470 data_array.data0\[4\]\[2\] VGND VGND VPWR VPWR net2121 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold481 tag_array.tag1\[2\]\[17\] VGND VGND VPWR VPWR net2132 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold492 data_array.data0\[2\]\[15\] VGND VGND VPWR VPWR net2143 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_225_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_225_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11011_ net2532 net956 net341 VGND VGND VPWR VPWR _02755_ sky130_fd_sc_hd__mux2_1
Xfanout950 _05500_ VGND VGND VPWR VPWR net950 sky130_fd_sc_hd__clkbuf_2
Xfanout961 net963 VGND VGND VPWR VPWR net961 sky130_fd_sc_hd__clkbuf_2
XFILLER_131_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout972 _05488_ VGND VGND VPWR VPWR net972 sky130_fd_sc_hd__clkbuf_2
Xfanout983 _05484_ VGND VGND VPWR VPWR net983 sky130_fd_sc_hd__buf_1
XFILLER_86_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout994 net995 VGND VGND VPWR VPWR net994 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12962_ clknet_leaf_168_clk _01656_ VGND VGND VPWR VPWR tag_array.tag0\[4\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1170 data_array.data0\[5\]\[7\] VGND VGND VPWR VPWR net2821 sky130_fd_sc_hd__dlygate4sd3_1
X_11913_ clknet_leaf_1_clk _00721_ VGND VGND VPWR VPWR data_array.data0\[5\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1181 data_array.data1\[6\]\[37\] VGND VGND VPWR VPWR net2832 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1192 tag_array.tag0\[12\]\[20\] VGND VGND VPWR VPWR net2843 sky130_fd_sc_hd__dlygate4sd3_1
X_12893_ clknet_leaf_205_clk _01587_ VGND VGND VPWR VPWR data_array.data0\[12\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_46_878 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11844_ clknet_leaf_243_clk _00652_ VGND VGND VPWR VPWR data_array.data0\[7\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_68_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11775_ clknet_leaf_259_clk _00583_ VGND VGND VPWR VPWR data_array.data0\[8\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10726_ net1070 net2761 net500 VGND VGND VPWR VPWR _02471_ sky130_fd_sc_hd__mux2_1
X_13514_ clknet_leaf_35_clk _02143_ VGND VGND VPWR VPWR data_array.data1\[0\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14494_ clknet_leaf_162_clk _03117_ VGND VGND VPWR VPWR tag_array.dirty0\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_13_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13445_ clknet_leaf_166_clk _02075_ VGND VGND VPWR VPWR tag_array.tag0\[1\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_146_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10657_ net2071 net1090 net482 VGND VGND VPWR VPWR _02402_ sky130_fd_sc_hd__mux2_1
XFILLER_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload15 clknet_leaf_0_clk VGND VGND VPWR VPWR clkload15/Y sky130_fd_sc_hd__inv_6
Xclkload26 clknet_leaf_265_clk VGND VGND VPWR VPWR clkload26/Y sky130_fd_sc_hd__inv_8
XFILLER_10_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload37 clknet_leaf_7_clk VGND VGND VPWR VPWR clkload37/Y sky130_fd_sc_hd__clkinv_8
XFILLER_62_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13376_ clknet_leaf_162_clk _02006_ VGND VGND VPWR VPWR tag_array.tag0\[2\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_10588_ net2581 net1110 net477 VGND VGND VPWR VPWR _02333_ sky130_fd_sc_hd__mux2_1
XFILLER_182_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload48 clknet_leaf_258_clk VGND VGND VPWR VPWR clkload48/Y sky130_fd_sc_hd__clkinv_2
XFILLER_5_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload59 clknet_leaf_25_clk VGND VGND VPWR VPWR clkload59/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_115_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12327_ clknet_leaf_62_clk _00063_ VGND VGND VPWR VPWR data_array.rdata0\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_142_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12258_ clknet_leaf_98_clk _01016_ VGND VGND VPWR VPWR tag_array.tag1\[14\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_216_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_216_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_68_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11209_ net937 net3204 net655 VGND VGND VPWR VPWR _02952_ sky130_fd_sc_hd__mux2_1
X_12189_ clknet_leaf_155_clk _00997_ VGND VGND VPWR VPWR tag_array.tag0\[14\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_110_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1032 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06750_ data_array.data0\[1\]\[1\] net1523 net1427 data_array.data0\[2\]\[1\] VGND
+ VGND VPWR VPWR _04054_ sky130_fd_sc_hd__a22o_1
XFILLER_83_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_108_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05701_ fsm.tag_out0\[1\] net31 VGND VGND VPWR VPWR _03218_ sky130_fd_sc_hd__and2b_1
X_06681_ _03990_ _03991_ VGND VGND VPWR VPWR _00166_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_125_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08420_ net1884 net916 net692 VGND VGND VPWR VPWR _00269_ sky130_fd_sc_hd__mux2_1
XFILLER_52_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05632_ _03150_ VGND VGND VPWR VPWR _03151_ sky130_fd_sc_hd__inv_2
XFILLER_52_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08351_ net2424 net1010 net686 VGND VGND VPWR VPWR _00246_ sky130_fd_sc_hd__mux2_1
XFILLER_177_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07302_ data_array.data0\[9\]\[51\] net1522 net1426 data_array.data0\[10\]\[51\]
+ VGND VGND VPWR VPWR _04556_ sky130_fd_sc_hd__a22o_1
XFILLER_20_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08282_ net2043 net1102 net689 VGND VGND VPWR VPWR _00223_ sky130_fd_sc_hd__mux2_1
XFILLER_149_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload9 clknet_5_20__leaf_clk VGND VGND VPWR VPWR clkload9/X sky130_fd_sc_hd__clkbuf_8
X_07233_ data_array.data0\[12\]\[45\] net1344 net1250 data_array.data0\[15\]\[45\]
+ _04492_ VGND VGND VPWR VPWR _04493_ sky130_fd_sc_hd__a221o_1
XFILLER_177_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07164_ net1227 _04425_ _04429_ net1179 VGND VGND VPWR VPWR _04431_ sky130_fd_sc_hd__a22o_1
XFILLER_145_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06115_ data_array.rdata0\[30\] net1139 net1115 data_array.rdata1\[30\] VGND VGND
+ VPWR VPWR net286 sky130_fd_sc_hd__a22o_1
XFILLER_117_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07095_ data_array.data0\[5\]\[32\] net1520 net1424 data_array.data0\[6\]\[32\] VGND
+ VGND VPWR VPWR _04368_ sky130_fd_sc_hd__a22o_1
XFILLER_118_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06046_ net1653 net1121 _03486_ VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__a21o_1
XFILLER_160_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_207_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_207_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_132_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_184_3887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_184_3898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09805_ net988 net3367 net391 VGND VGND VPWR VPWR _01556_ sky130_fd_sc_hd__mux2_1
X_07997_ data_array.data1\[1\]\[50\] net1527 net1431 data_array.data1\[2\]\[50\] VGND
+ VGND VPWR VPWR _05188_ sky130_fd_sc_hd__a22o_1
XFILLER_75_17 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06948_ data_array.data0\[5\]\[19\] net1581 net1485 data_array.data0\[6\]\[19\] VGND
+ VGND VPWR VPWR _04234_ sky130_fd_sc_hd__a22o_1
X_09736_ net742 net3953 net679 VGND VGND VPWR VPWR _01488_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09667_ net720 net3664 net612 VGND VGND VPWR VPWR _01419_ sky130_fd_sc_hd__mux2_1
X_06879_ _04170_ _04171_ VGND VGND VPWR VPWR _00003_ sky130_fd_sc_hd__or2_1
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08618_ net750 net2613 net523 VGND VGND VPWR VPWR _00377_ sky130_fd_sc_hd__mux2_1
X_09598_ net957 net3874 net398 VGND VGND VPWR VPWR _01350_ sky130_fd_sc_hd__mux2_1
XFILLER_70_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08549_ net760 net2653 net589 VGND VGND VPWR VPWR _00317_ sky130_fd_sc_hd__mux2_1
XFILLER_39_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11560_ clknet_leaf_32_clk _00368_ VGND VGND VPWR VPWR tag_array.tag1\[5\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_168_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10511_ net903 net2944 net346 VGND VGND VPWR VPWR _02256_ sky130_fd_sc_hd__mux2_1
XFILLER_7_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11491_ clknet_leaf_153_clk _00300_ VGND VGND VPWR VPWR tag_array.valid0\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_11_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13230_ clknet_leaf_47_clk _01860_ VGND VGND VPWR VPWR data_array.data0\[11\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_137_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10442_ net2051 net886 net663 VGND VGND VPWR VPWR _02188_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_21_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13161_ clknet_leaf_130_clk _01855_ VGND VGND VPWR VPWR tag_array.tag1\[8\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_152_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10373_ net708 net2879 net539 VGND VGND VPWR VPWR _02120_ sky130_fd_sc_hd__mux2_1
XFILLER_151_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12112_ clknet_leaf_203_clk _00920_ VGND VGND VPWR VPWR data_array.data1\[14\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_163_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13092_ clknet_leaf_43_clk _01786_ VGND VGND VPWR VPWR data_array.data1\[13\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_151_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12043_ clknet_leaf_2_clk _00851_ VGND VGND VPWR VPWR data_array.data0\[6\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_133_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout780 net781 VGND VGND VPWR VPWR net780 sky130_fd_sc_hd__buf_1
XFILLER_37_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout791 net792 VGND VGND VPWR VPWR net791 sky130_fd_sc_hd__clkbuf_2
X_13994_ clknet_leaf_8_clk _02623_ VGND VGND VPWR VPWR data_array.data1\[5\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12945_ clknet_leaf_53_clk _01639_ VGND VGND VPWR VPWR data_array.data0\[13\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_142_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12876_ clknet_leaf_84_clk _01570_ VGND VGND VPWR VPWR data_array.data0\[12\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11827_ clknet_leaf_52_clk _00635_ VGND VGND VPWR VPWR data_array.data0\[7\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_83_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_120_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11758_ clknet_leaf_96_clk _00566_ VGND VGND VPWR VPWR data_array.data0\[8\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_10709_ net2403 net883 net478 VGND VGND VPWR VPWR _02454_ sky130_fd_sc_hd__mux2_1
X_11689_ clknet_leaf_136_clk _00497_ VGND VGND VPWR VPWR tag_array.tag1\[15\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_14477_ clknet_leaf_211_clk _03100_ VGND VGND VPWR VPWR data_array.data1\[7\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload104 clknet_leaf_39_clk VGND VGND VPWR VPWR clkload104/X sky130_fd_sc_hd__clkbuf_8
X_13428_ clknet_leaf_76_clk _02058_ VGND VGND VPWR VPWR data_array.data1\[8\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload115 clknet_leaf_98_clk VGND VGND VPWR VPWR clkload115/Y sky130_fd_sc_hd__clkinv_4
XFILLER_139_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload126 clknet_leaf_81_clk VGND VGND VPWR VPWR clkload126/Y sky130_fd_sc_hd__inv_8
Xclkload137 clknet_leaf_219_clk VGND VGND VPWR VPWR clkload137/Y sky130_fd_sc_hd__inv_8
Xclkload148 clknet_leaf_225_clk VGND VGND VPWR VPWR clkload148/Y sky130_fd_sc_hd__inv_6
Xclkload159 clknet_leaf_172_clk VGND VGND VPWR VPWR clkload159/Y sky130_fd_sc_hd__clkinvlp_4
X_13359_ clknet_leaf_191_clk _01989_ VGND VGND VPWR VPWR tag_array.tag0\[2\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_149_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_149_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07920_ data_array.data1\[5\]\[43\] net1568 net1472 data_array.data1\[6\]\[43\] VGND
+ VGND VPWR VPWR _05118_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_166_3551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2607 data_array.data1\[10\]\[32\] VGND VGND VPWR VPWR net4258 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2618 data_array.data0\[3\]\[38\] VGND VGND VPWR VPWR net4269 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2629 data_array.data1\[4\]\[35\] VGND VGND VPWR VPWR net4280 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07851_ data_array.data1\[0\]\[37\] net1353 net1259 data_array.data1\[3\]\[37\] _05054_
+ VGND VGND VPWR VPWR _05055_ sky130_fd_sc_hd__a221o_1
Xhold1906 data_array.data1\[14\]\[43\] VGND VGND VPWR VPWR net3557 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_127_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1917 data_array.data1\[12\]\[24\] VGND VGND VPWR VPWR net3568 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1928 data_array.data1\[3\]\[21\] VGND VGND VPWR VPWR net3579 sky130_fd_sc_hd__dlygate4sd3_1
X_06802_ _04100_ _04101_ VGND VGND VPWR VPWR _00055_ sky130_fd_sc_hd__or2_1
Xhold1939 data_array.data1\[6\]\[2\] VGND VGND VPWR VPWR net3590 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput2 cpu_addr[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_2
X_07782_ data_array.data1\[13\]\[31\] net1576 net1480 data_array.data1\[14\]\[31\]
+ VGND VGND VPWR VPWR _04992_ sky130_fd_sc_hd__a22o_1
XFILLER_68_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09521_ net745 net2106 net621 VGND VGND VPWR VPWR _01274_ sky130_fd_sc_hd__mux2_1
X_06733_ tag_array.tag1\[0\]\[24\] net1372 net1278 tag_array.tag1\[3\]\[24\] _04038_
+ VGND VGND VPWR VPWR _04039_ sky130_fd_sc_hd__a221o_1
XFILLER_37_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09452_ net859 net2545 net583 VGND VGND VPWR VPWR _01205_ sky130_fd_sc_hd__mux2_1
XFILLER_52_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06664_ tag_array.tag1\[9\]\[18\] net1562 net1466 tag_array.tag1\[10\]\[18\] VGND
+ VGND VPWR VPWR _03976_ sky130_fd_sc_hd__a22o_1
XFILLER_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08403_ net136 net71 net1640 VGND VGND VPWR VPWR _05505_ sky130_fd_sc_hd__mux2_1
XFILLER_149_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05615_ fsm.tag_out1\[3\] VGND VGND VPWR VPWR _03137_ sky130_fd_sc_hd__inv_2
X_09383_ net868 net2999 net408 VGND VGND VPWR VPWR _01136_ sky130_fd_sc_hd__mux2_1
XFILLER_80_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06595_ tag_array.tag1\[12\]\[12\] net1401 net1307 tag_array.tag1\[15\]\[12\] _03912_
+ VGND VGND VPWR VPWR _03913_ sky130_fd_sc_hd__a221o_1
X_08334_ net111 net46 net1648 VGND VGND VPWR VPWR _05459_ sky130_fd_sc_hd__mux2_1
XFILLER_20_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08265_ net700 net4116 net805 VGND VGND VPWR VPWR _00219_ sky130_fd_sc_hd__mux2_1
X_07216_ data_array.data0\[5\]\[43\] net1567 net1471 data_array.data0\[6\]\[43\] VGND
+ VGND VPWR VPWR _04478_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_41_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08196_ net791 net3518 net800 VGND VGND VPWR VPWR _00196_ sky130_fd_sc_hd__mux2_1
X_07147_ data_array.data0\[0\]\[37\] net1353 net1259 data_array.data0\[3\]\[37\] _04414_
+ VGND VGND VPWR VPWR _04415_ sky130_fd_sc_hd__a221o_1
XFILLER_134_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_1013 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07078_ data_array.data0\[13\]\[31\] net1574 net1478 data_array.data0\[14\]\[31\]
+ VGND VGND VPWR VPWR _04352_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_7_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06029_ fsm.lru_out fsm.valid1 fsm.state\[5\] VGND VGND VPWR VPWR _03479_ sky130_fd_sc_hd__and3_1
XFILLER_126_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1008 net1011 VGND VGND VPWR VPWR net1008 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1019 _05466_ VGND VGND VPWR VPWR net1019 sky130_fd_sc_hd__buf_1
XFILLER_114_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09719_ net712 net2467 net609 VGND VGND VPWR VPWR _01471_ sky130_fd_sc_hd__mux2_1
XFILLER_74_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10991_ net2368 net1036 net337 VGND VGND VPWR VPWR _02735_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12730_ clknet_leaf_108_clk _01424_ VGND VGND VPWR VPWR tag_array.tag0\[7\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12661_ clknet_leaf_47_clk _01355_ VGND VGND VPWR VPWR data_array.data0\[15\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_26_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11612_ clknet_leaf_191_clk _00420_ VGND VGND VPWR VPWR tag_array.tag1\[3\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_14400_ clknet_leaf_242_clk _03023_ VGND VGND VPWR VPWR data_array.data1\[10\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_26_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12592_ clknet_leaf_185_clk _01286_ VGND VGND VPWR VPWR tag_array.tag0\[10\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_5_19__f_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_5_19__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_61_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14331_ clknet_leaf_5_clk _02960_ VGND VGND VPWR VPWR data_array.data1\[11\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
X_11543_ clknet_leaf_127_clk _00351_ VGND VGND VPWR VPWR tag_array.tag1\[6\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14262_ clknet_leaf_6_clk _02891_ VGND VGND VPWR VPWR data_array.data1\[12\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
X_11474_ clknet_leaf_224_clk _00284_ VGND VGND VPWR VPWR data_array.data0\[0\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13213_ clknet_leaf_253_clk _00109_ VGND VGND VPWR VPWR data_array.rdata1\[50\] sky130_fd_sc_hd__dfxtp_1
X_10425_ net2164 net952 net663 VGND VGND VPWR VPWR _02171_ sky130_fd_sc_hd__mux2_1
XFILLER_137_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14193_ clknet_leaf_260_clk _02822_ VGND VGND VPWR VPWR data_array.data0\[2\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_100_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13144_ clknet_leaf_195_clk _01838_ VGND VGND VPWR VPWR tag_array.tag1\[8\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_10356_ net776 net4392 net538 VGND VGND VPWR VPWR _02103_ sky130_fd_sc_hd__mux2_1
XFILLER_100_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13075_ clknet_leaf_255_clk _01769_ VGND VGND VPWR VPWR data_array.data1\[13\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_10287_ net2241 net1014 net641 VGND VGND VPWR VPWR _02034_ sky130_fd_sc_hd__mux2_1
X_12026_ clknet_leaf_113_clk _00834_ VGND VGND VPWR VPWR data_array.data0\[6\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout1520 net1521 VGND VGND VPWR VPWR net1520 sky130_fd_sc_hd__clkbuf_4
Xfanout1531 net1533 VGND VGND VPWR VPWR net1531 sky130_fd_sc_hd__clkbuf_4
Xfanout1542 net1543 VGND VGND VPWR VPWR net1542 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_144_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1553 net1554 VGND VGND VPWR VPWR net1553 sky130_fd_sc_hd__clkbuf_4
Xfanout1564 net1565 VGND VGND VPWR VPWR net1564 sky130_fd_sc_hd__clkbuf_4
Xfanout1575 net1576 VGND VGND VPWR VPWR net1575 sky130_fd_sc_hd__clkbuf_4
XFILLER_65_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1586 net1587 VGND VGND VPWR VPWR net1586 sky130_fd_sc_hd__clkbuf_4
XFILLER_76_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1597 net1600 VGND VGND VPWR VPWR net1597 sky130_fd_sc_hd__clkbuf_4
XFILLER_53_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13977_ clknet_leaf_254_clk _02606_ VGND VGND VPWR VPWR data_array.data1\[5\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_122_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12928_ clknet_leaf_261_clk _01622_ VGND VGND VPWR VPWR data_array.data0\[13\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_179_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12859_ clknet_leaf_237_clk _01553_ VGND VGND VPWR VPWR data_array.data0\[12\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_06380_ tag_array.tag0\[1\]\[17\] net1602 net1506 tag_array.tag0\[2\]\[17\] VGND
+ VGND VPWR VPWR _03718_ sky130_fd_sc_hd__a22o_1
XFILLER_175_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_1_Left_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08050_ data_array.data1\[9\]\[55\] net1535 net1439 data_array.data1\[10\]\[55\]
+ VGND VGND VPWR VPWR _05236_ sky130_fd_sc_hd__a22o_1
XFILLER_179_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07001_ data_array.data0\[13\]\[24\] net1575 net1479 data_array.data0\[14\]\[24\]
+ VGND VGND VPWR VPWR _04282_ sky130_fd_sc_hd__a22o_1
XFILLER_115_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08952_ net956 net4155 net430 VGND VGND VPWR VPWR _00708_ sky130_fd_sc_hd__mux2_1
XFILLER_115_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2404 data_array.data0\[11\]\[21\] VGND VGND VPWR VPWR net4055 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2415 data_array.data0\[13\]\[52\] VGND VGND VPWR VPWR net4066 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_181_3835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07903_ data_array.data1\[9\]\[42\] net1585 net1489 data_array.data1\[10\]\[42\]
+ VGND VGND VPWR VPWR _05102_ sky130_fd_sc_hd__a22o_1
Xhold2426 data_array.data1\[14\]\[51\] VGND VGND VPWR VPWR net4077 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_181_3846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08883_ net972 net4114 net435 VGND VGND VPWR VPWR _00640_ sky130_fd_sc_hd__mux2_1
Xhold2437 data_array.data0\[10\]\[50\] VGND VGND VPWR VPWR net4088 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2448 tag_array.tag1\[15\]\[14\] VGND VGND VPWR VPWR net4099 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1703 data_array.data0\[9\]\[48\] VGND VGND VPWR VPWR net3354 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1714 data_array.data1\[10\]\[38\] VGND VGND VPWR VPWR net3365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2459 data_array.data1\[14\]\[2\] VGND VGND VPWR VPWR net4110 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1725 data_array.data0\[15\]\[18\] VGND VGND VPWR VPWR net3376 sky130_fd_sc_hd__dlygate4sd3_1
X_07834_ net1190 _05033_ _05037_ net1616 VGND VGND VPWR VPWR _05040_ sky130_fd_sc_hd__a22o_1
XFILLER_57_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1736 tag_array.tag1\[6\]\[15\] VGND VGND VPWR VPWR net3387 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1747 data_array.data1\[14\]\[21\] VGND VGND VPWR VPWR net3398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1758 data_array.data1\[7\]\[19\] VGND VGND VPWR VPWR net3409 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_99_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_556 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1769 tag_array.tag0\[6\]\[2\] VGND VGND VPWR VPWR net3420 sky130_fd_sc_hd__dlygate4sd3_1
X_07765_ data_array.data1\[8\]\[29\] net1387 net1293 data_array.data1\[11\]\[29\]
+ _04976_ VGND VGND VPWR VPWR _04977_ sky130_fd_sc_hd__a221o_1
XFILLER_84_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06716_ tag_array.tag1\[8\]\[23\] net1419 net1325 tag_array.tag1\[11\]\[23\] _04022_
+ VGND VGND VPWR VPWR _04023_ sky130_fd_sc_hd__a221o_1
XFILLER_65_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09504_ net712 net2775 net624 VGND VGND VPWR VPWR _01257_ sky130_fd_sc_hd__mux2_1
X_07696_ data_array.data1\[1\]\[23\] net1550 net1454 data_array.data1\[2\]\[23\] VGND
+ VGND VPWR VPWR _04914_ sky130_fd_sc_hd__a22o_1
XFILLER_112_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09435_ net924 net2770 net578 VGND VGND VPWR VPWR _01188_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_179_3797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06647_ net1232 _03955_ _03959_ net1184 VGND VGND VPWR VPWR _03961_ sky130_fd_sc_hd__a22o_1
XFILLER_52_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09366_ net936 net4414 net406 VGND VGND VPWR VPWR _01119_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06578_ tag_array.tag1\[5\]\[10\] net1596 net1500 tag_array.tag1\[6\]\[10\] VGND
+ VGND VPWR VPWR _03898_ sky130_fd_sc_hd__a22o_1
X_08317_ net1128 _05447_ VGND VGND VPWR VPWR _05448_ sky130_fd_sc_hd__and2_1
XANTENNA_40 net493 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09297_ net792 net2516 net548 VGND VGND VPWR VPWR _01051_ sky130_fd_sc_hd__mux2_1
XANTENNA_51 net1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_62 net1518 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_73 _03153_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08248_ _03142_ _03147_ VGND VGND VPWR VPWR _05400_ sky130_fd_sc_hd__nor2_1
XANTENNA_84 net1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_826 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08179_ net849 _03285_ net4614 VGND VGND VPWR VPWR _00183_ sky130_fd_sc_hd__a21boi_1
X_10210_ net965 net2768 net360 VGND VGND VPWR VPWR _01957_ sky130_fd_sc_hd__mux2_1
XFILLER_118_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_904 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11190_ net1014 net3312 net656 VGND VGND VPWR VPWR _02933_ sky130_fd_sc_hd__mux2_1
XFILLER_134_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10141_ net983 net4498 net362 VGND VGND VPWR VPWR _01889_ sky130_fd_sc_hd__mux2_1
Xoutput180 net180 VGND VGND VPWR VPWR cpu_rdata[23] sky130_fd_sc_hd__clkbuf_4
Xoutput191 net191 VGND VGND VPWR VPWR cpu_rdata[33] sky130_fd_sc_hd__buf_6
XFILLER_82_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10072_ net735 net3840 net599 VGND VGND VPWR VPWR _01821_ sky130_fd_sc_hd__mux2_1
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13900_ clknet_leaf_69_clk _02529_ VGND VGND VPWR VPWR data_array.data1\[4\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2960 data_array.data1\[13\]\[39\] VGND VGND VPWR VPWR net4611 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2971 tag_array.tag1\[5\]\[9\] VGND VGND VPWR VPWR net4622 sky130_fd_sc_hd__dlygate4sd3_1
X_13831_ clknet_leaf_192_clk _02460_ VGND VGND VPWR VPWR data_array.data1\[2\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10974_ net3039 net1105 net336 VGND VGND VPWR VPWR _02718_ sky130_fd_sc_hd__mux2_1
X_13762_ clknet_leaf_202_clk _02391_ VGND VGND VPWR VPWR data_array.data1\[1\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12713_ clknet_leaf_181_clk _01407_ VGND VGND VPWR VPWR tag_array.tag0\[7\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_100_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13693_ clknet_leaf_5_clk _02322_ VGND VGND VPWR VPWR data_array.data1\[15\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_80_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12644_ clknet_leaf_245_clk _01338_ VGND VGND VPWR VPWR data_array.data0\[15\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_129_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12575_ clknet_leaf_143_clk _01269_ VGND VGND VPWR VPWR tag_array.tag0\[10\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_873 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14314_ clknet_leaf_6_clk _02943_ VGND VGND VPWR VPWR data_array.data1\[11\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_157_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11526_ clknet_leaf_174_clk _00334_ VGND VGND VPWR VPWR tag_array.valid1\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_184_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11457_ clknet_leaf_23_clk _00267_ VGND VGND VPWR VPWR data_array.data0\[0\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
X_14245_ clknet_leaf_39_clk _02874_ VGND VGND VPWR VPWR data_array.data1\[12\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_171_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10408_ net2787 net1021 net663 VGND VGND VPWR VPWR _02154_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14176_ clknet_leaf_92_clk _02805_ VGND VGND VPWR VPWR data_array.data0\[2\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_11388_ clknet_leaf_233_clk _00198_ VGND VGND VPWR VPWR tag_array.tag1\[7\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_115_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_712 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13127_ clknet_leaf_231_clk _01821_ VGND VGND VPWR VPWR tag_array.tag0\[3\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_10339_ net745 net3055 net591 VGND VGND VPWR VPWR _02086_ sky130_fd_sc_hd__mux2_1
XFILLER_97_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_111_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ clknet_leaf_57_clk _01752_ VGND VGND VPWR VPWR data_array.data1\[13\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_140_778 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1350 net1352 VGND VGND VPWR VPWR net1350 sky130_fd_sc_hd__clkbuf_4
X_12009_ clknet_leaf_58_clk _00817_ VGND VGND VPWR VPWR data_array.data0\[6\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout1361 net1363 VGND VGND VPWR VPWR net1361 sky130_fd_sc_hd__clkbuf_4
X_05880_ data_array.rdata1\[16\] net830 net839 VGND VGND VPWR VPWR _03381_ sky130_fd_sc_hd__a21o_1
XFILLER_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1372 net1375 VGND VGND VPWR VPWR net1372 sky130_fd_sc_hd__clkbuf_4
Xfanout1383 net1400 VGND VGND VPWR VPWR net1383 sky130_fd_sc_hd__clkbuf_2
Xfanout1394 net1400 VGND VGND VPWR VPWR net1394 sky130_fd_sc_hd__clkbuf_4
XFILLER_38_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07550_ _04780_ _04781_ VGND VGND VPWR VPWR _00127_ sky130_fd_sc_hd__or2_1
XFILLER_19_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06501_ tag_array.tag1\[1\]\[3\] net1561 net1465 tag_array.tag1\[2\]\[3\] VGND VGND
+ VPWR VPWR _03828_ sky130_fd_sc_hd__a22o_1
X_07481_ data_array.data1\[0\]\[3\] net1384 net1290 data_array.data1\[3\]\[3\] _04718_
+ VGND VGND VPWR VPWR _04719_ sky130_fd_sc_hd__a221o_1
XFILLER_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09220_ net698 net2668 net631 VGND VGND VPWR VPWR _00974_ sky130_fd_sc_hd__mux2_1
X_06432_ tag_array.tag0\[4\]\[22\] net1374 net1280 tag_array.tag0\[7\]\[22\] _03764_
+ VGND VGND VPWR VPWR _03765_ sky130_fd_sc_hd__a221o_1
XFILLER_107_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09151_ net938 net3557 net573 VGND VGND VPWR VPWR _00905_ sky130_fd_sc_hd__mux2_1
X_06363_ tag_array.tag0\[9\]\[16\] net1598 net1502 tag_array.tag0\[10\]\[16\] VGND
+ VGND VPWR VPWR _03702_ sky130_fd_sc_hd__a22o_1
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08102_ data_array.data1\[8\]\[60\] net1414 net1320 data_array.data1\[11\]\[60\]
+ _05282_ VGND VGND VPWR VPWR _05283_ sky130_fd_sc_hd__a221o_1
XFILLER_30_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09082_ net956 net3341 net414 VGND VGND VPWR VPWR _00836_ sky130_fd_sc_hd__mux2_1
XFILLER_174_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06294_ net1208 _03633_ _03637_ net1634 VGND VGND VPWR VPWR _03640_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_135_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08033_ net1213 _05215_ _05219_ net1165 VGND VGND VPWR VPWR _05221_ sky130_fd_sc_hd__a22o_1
Xinput60 cpu_wdata[33] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_1
Xhold800 tag_array.tag0\[13\]\[0\] VGND VGND VPWR VPWR net2451 sky130_fd_sc_hd__dlygate4sd3_1
Xhold811 data_array.data0\[14\]\[19\] VGND VGND VPWR VPWR net2462 sky130_fd_sc_hd__dlygate4sd3_1
Xinput71 cpu_wdata[43] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_1
Xinput82 cpu_wdata[53] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_1
Xhold822 data_array.data0\[5\]\[19\] VGND VGND VPWR VPWR net2473 sky130_fd_sc_hd__dlygate4sd3_1
Xinput93 cpu_wdata[63] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_1
Xhold833 data_array.data1\[0\]\[52\] VGND VGND VPWR VPWR net2484 sky130_fd_sc_hd__dlygate4sd3_1
Xhold844 data_array.data0\[11\]\[48\] VGND VGND VPWR VPWR net2495 sky130_fd_sc_hd__dlygate4sd3_1
Xhold855 data_array.data1\[11\]\[5\] VGND VGND VPWR VPWR net2506 sky130_fd_sc_hd__dlygate4sd3_1
Xhold866 tag_array.tag1\[5\]\[18\] VGND VGND VPWR VPWR net2517 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold877 tag_array.tag1\[2\]\[7\] VGND VGND VPWR VPWR net2528 sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 tag_array.tag0\[12\]\[9\] VGND VGND VPWR VPWR net2539 sky130_fd_sc_hd__dlygate4sd3_1
Xhold899 data_array.data0\[1\]\[2\] VGND VGND VPWR VPWR net2550 sky130_fd_sc_hd__dlygate4sd3_1
X_09984_ net894 net4427 net372 VGND VGND VPWR VPWR _01733_ sky130_fd_sc_hd__mux2_1
XFILLER_107_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2201 data_array.data1\[9\]\[52\] VGND VGND VPWR VPWR net3852 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2212 tag_array.tag1\[14\]\[23\] VGND VGND VPWR VPWR net3863 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_67_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2223 data_array.data0\[15\]\[38\] VGND VGND VPWR VPWR net3874 sky130_fd_sc_hd__dlygate4sd3_1
X_08935_ net1025 net4473 net428 VGND VGND VPWR VPWR _00691_ sky130_fd_sc_hd__mux2_1
XFILLER_76_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2234 data_array.data0\[15\]\[55\] VGND VGND VPWR VPWR net3885 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_36_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2245 data_array.data0\[7\]\[12\] VGND VGND VPWR VPWR net3896 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1500 data_array.data0\[5\]\[42\] VGND VGND VPWR VPWR net3151 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1511 data_array.data0\[7\]\[41\] VGND VGND VPWR VPWR net3162 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2256 data_array.data0\[3\]\[47\] VGND VGND VPWR VPWR net3907 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2267 tag_array.dirty1\[12\] VGND VGND VPWR VPWR net3918 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1522 tag_array.tag1\[15\]\[10\] VGND VGND VPWR VPWR net3173 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2278 data_array.data1\[13\]\[33\] VGND VGND VPWR VPWR net3929 sky130_fd_sc_hd__dlygate4sd3_1
X_08866_ net1042 net2461 net436 VGND VGND VPWR VPWR _00623_ sky130_fd_sc_hd__mux2_1
Xhold1533 data_array.data1\[2\]\[28\] VGND VGND VPWR VPWR net3184 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1544 tag_array.tag0\[12\]\[3\] VGND VGND VPWR VPWR net3195 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2289 tag_array.tag1\[6\]\[13\] VGND VGND VPWR VPWR net3940 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1555 data_array.data1\[10\]\[16\] VGND VGND VPWR VPWR net3206 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07817_ data_array.data1\[5\]\[34\] net1531 net1435 data_array.data1\[6\]\[34\] VGND
+ VGND VPWR VPWR _05024_ sky130_fd_sc_hd__a22o_1
XFILLER_84_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1566 data_array.data0\[9\]\[29\] VGND VGND VPWR VPWR net3217 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1577 tag_array.tag1\[15\]\[22\] VGND VGND VPWR VPWR net3228 sky130_fd_sc_hd__dlygate4sd3_1
X_08797_ net3325 net1059 net444 VGND VGND VPWR VPWR _00555_ sky130_fd_sc_hd__mux2_1
Xhold1588 data_array.data1\[13\]\[14\] VGND VGND VPWR VPWR net3239 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1599 data_array.data0\[3\]\[44\] VGND VGND VPWR VPWR net3250 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_28_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07748_ _04960_ _04961_ VGND VGND VPWR VPWR _00083_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_64_Left_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07679_ data_array.data1\[4\]\[21\] net1365 net1271 data_array.data1\[7\]\[21\] _04898_
+ VGND VGND VPWR VPWR _04899_ sky130_fd_sc_hd__a221o_1
XFILLER_13_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09418_ net994 net3736 net585 VGND VGND VPWR VPWR _01171_ sky130_fd_sc_hd__mux2_1
X_10690_ net2287 net957 net485 VGND VGND VPWR VPWR _02435_ sky130_fd_sc_hd__mux2_1
XFILLER_12_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09349_ net1006 net2958 net403 VGND VGND VPWR VPWR _01102_ sky130_fd_sc_hd__mux2_1
X_12360_ clknet_leaf_80_clk _00036_ VGND VGND VPWR VPWR data_array.rdata0\[42\] sky130_fd_sc_hd__dfxtp_1
X_11311_ net1051 net3488 net801 VGND VGND VPWR VPWR _03054_ sky130_fd_sc_hd__mux2_1
X_12291_ clknet_leaf_130_clk _01049_ VGND VGND VPWR VPWR tag_array.tag1\[13\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_180_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14030_ clknet_leaf_269_clk _02659_ VGND VGND VPWR VPWR data_array.data1\[6\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11242_ net1063 net4169 net682 VGND VGND VPWR VPWR _02985_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_73_Left_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11173_ net1082 net3069 net657 VGND VGND VPWR VPWR _02916_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10124_ net1049 net1894 net367 VGND VGND VPWR VPWR _01872_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_73_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10055_ net864 net2777 net558 VGND VGND VPWR VPWR _01804_ sky130_fd_sc_hd__mux2_1
XFILLER_180_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2790 data_array.data0\[11\]\[11\] VGND VGND VPWR VPWR net4441 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13814_ clknet_leaf_5_clk _02443_ VGND VGND VPWR VPWR data_array.data1\[2\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_82_Left_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13745_ clknet_leaf_257_clk _02374_ VGND VGND VPWR VPWR data_array.data1\[1\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
X_10957_ net915 net4086 net532 VGND VGND VPWR VPWR _02702_ sky130_fd_sc_hd__mux2_1
XFILLER_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13676_ clknet_leaf_118_clk _02305_ VGND VGND VPWR VPWR data_array.data1\[15\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
X_10888_ net934 net2665 net521 VGND VGND VPWR VPWR _02633_ sky130_fd_sc_hd__mux2_1
XFILLER_176_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12627_ clknet_leaf_61_clk _01321_ VGND VGND VPWR VPWR data_array.data0\[15\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12558_ clknet_leaf_162_clk _01252_ VGND VGND VPWR VPWR tag_array.tag0\[11\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_152_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11509_ clknet_leaf_137_clk _00317_ VGND VGND VPWR VPWR tag_array.tag1\[9\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_91_Left_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12489_ clknet_leaf_260_clk _01183_ VGND VGND VPWR VPWR data_array.data1\[9\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold107 tag_array.tag1\[1\]\[15\] VGND VGND VPWR VPWR net1758 sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 data_array.data1\[0\]\[31\] VGND VGND VPWR VPWR net1769 sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 data_array.data1\[2\]\[2\] VGND VGND VPWR VPWR net1780 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14228_ clknet_leaf_85_clk _02857_ VGND VGND VPWR VPWR data_array.data1\[12\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_113_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14159_ clknet_leaf_113_clk _02788_ VGND VGND VPWR VPWR data_array.data0\[2\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout609 net611 VGND VGND VPWR VPWR net609 sky130_fd_sc_hd__buf_4
XFILLER_98_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06981_ data_array.data0\[1\]\[22\] net1532 net1436 data_array.data0\[2\]\[22\] VGND
+ VGND VPWR VPWR _04264_ sky130_fd_sc_hd__a22o_1
XFILLER_112_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05932_ net125 net1155 _03414_ _03415_ VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__a22o_1
X_08720_ net2917 net742 net476 VGND VGND VPWR VPWR _00479_ sky130_fd_sc_hd__mux2_1
XFILLER_78_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1180 net1187 VGND VGND VPWR VPWR net1180 sky130_fd_sc_hd__buf_4
Xfanout1191 net1212 VGND VGND VPWR VPWR net1191 sky130_fd_sc_hd__buf_2
X_08651_ net1827 net719 net513 VGND VGND VPWR VPWR _00410_ sky130_fd_sc_hd__mux2_1
X_05863_ net100 net1157 _03368_ _03369_ VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__a22o_1
XFILLER_82_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07602_ data_array.data1\[0\]\[14\] net1377 net1283 data_array.data1\[3\]\[14\] _04828_
+ VGND VGND VPWR VPWR _04829_ sky130_fd_sc_hd__a221o_1
X_08582_ net1721 net452 VGND VGND VPWR VPWR _00341_ sky130_fd_sc_hd__nand2b_1
XFILLER_81_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05794_ _03140_ fsm.tag_out1\[14\] _03243_ VGND VGND VPWR VPWR _03311_ sky130_fd_sc_hd__o21ai_1
XFILLER_183_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07533_ data_array.data1\[9\]\[8\] net1535 net1439 data_array.data1\[10\]\[8\] VGND
+ VGND VPWR VPWR _04766_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_176_3734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_176_3745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07464_ data_array.data1\[12\]\[2\] net1339 net1245 data_array.data1\[15\]\[2\] _04702_
+ VGND VGND VPWR VPWR _04703_ sky130_fd_sc_hd__a221o_1
XFILLER_22_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06415_ net1199 _03743_ _03747_ net1625 VGND VGND VPWR VPWR _03750_ sky130_fd_sc_hd__a22o_1
X_09203_ net769 net2996 net632 VGND VGND VPWR VPWR _00957_ sky130_fd_sc_hd__mux2_1
X_07395_ net1224 _04635_ _04639_ net1176 VGND VGND VPWR VPWR _04641_ sky130_fd_sc_hd__a22o_1
X_09134_ net1004 net3187 net567 VGND VGND VPWR VPWR _00888_ sky130_fd_sc_hd__mux2_1
X_06346_ tag_array.tag0\[12\]\[14\] net1369 net1275 tag_array.tag0\[15\]\[14\] _03686_
+ VGND VGND VPWR VPWR _03687_ sky130_fd_sc_hd__a221o_1
XFILLER_176_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09065_ net1025 net3955 net412 VGND VGND VPWR VPWR _00819_ sky130_fd_sc_hd__mux2_1
X_06277_ tag_array.tag0\[1\]\[8\] net1599 net1503 tag_array.tag0\[2\]\[8\] VGND VGND
+ VPWR VPWR _03624_ sky130_fd_sc_hd__a22o_1
XFILLER_162_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08016_ data_array.data1\[4\]\[52\] net1354 net1260 data_array.data1\[7\]\[52\] _05204_
+ VGND VGND VPWR VPWR _05205_ sky130_fd_sc_hd__a221o_1
Xhold630 data_array.data1\[1\]\[46\] VGND VGND VPWR VPWR net2281 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold641 data_array.data1\[4\]\[52\] VGND VGND VPWR VPWR net2292 sky130_fd_sc_hd__dlygate4sd3_1
Xhold652 data_array.data0\[1\]\[23\] VGND VGND VPWR VPWR net2303 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold663 tag_array.tag1\[11\]\[8\] VGND VGND VPWR VPWR net2314 sky130_fd_sc_hd__dlygate4sd3_1
Xhold674 data_array.data1\[1\]\[21\] VGND VGND VPWR VPWR net2325 sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 tag_array.tag1\[14\]\[17\] VGND VGND VPWR VPWR net2336 sky130_fd_sc_hd__dlygate4sd3_1
Xhold696 tag_array.tag1\[7\]\[5\] VGND VGND VPWR VPWR net2347 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_34_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09967_ net961 net2680 net372 VGND VGND VPWR VPWR _01716_ sky130_fd_sc_hd__mux2_1
XFILLER_58_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2020 data_array.data1\[11\]\[49\] VGND VGND VPWR VPWR net3671 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2031 data_array.data0\[11\]\[23\] VGND VGND VPWR VPWR net3682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2042 tag_array.tag1\[0\]\[9\] VGND VGND VPWR VPWR net3693 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2053 tag_array.tag1\[5\]\[4\] VGND VGND VPWR VPWR net3704 sky130_fd_sc_hd__dlygate4sd3_1
X_08918_ net1092 net3064 net431 VGND VGND VPWR VPWR _00674_ sky130_fd_sc_hd__mux2_1
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09898_ net877 net3443 net381 VGND VGND VPWR VPWR _01648_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_51_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2064 data_array.data1\[10\]\[3\] VGND VGND VPWR VPWR net3715 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2075 data_array.data1\[13\]\[28\] VGND VGND VPWR VPWR net3726 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1330 tag_array.tag0\[0\]\[8\] VGND VGND VPWR VPWR net2981 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1341 data_array.data0\[13\]\[8\] VGND VGND VPWR VPWR net2992 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2086 tag_array.tag0\[3\]\[12\] VGND VGND VPWR VPWR net3737 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1352 data_array.data0\[12\]\[32\] VGND VGND VPWR VPWR net3003 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2097 data_array.data1\[13\]\[6\] VGND VGND VPWR VPWR net3748 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1363 data_array.data1\[0\]\[6\] VGND VGND VPWR VPWR net3014 sky130_fd_sc_hd__dlygate4sd3_1
X_08849_ net1108 net3846 net437 VGND VGND VPWR VPWR _00606_ sky130_fd_sc_hd__mux2_1
XFILLER_85_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1374 data_array.data1\[14\]\[22\] VGND VGND VPWR VPWR net3025 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1385 data_array.data1\[13\]\[55\] VGND VGND VPWR VPWR net3036 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1396 tag_array.tag1\[13\]\[17\] VGND VGND VPWR VPWR net3047 sky130_fd_sc_hd__dlygate4sd3_1
X_11860_ clknet_leaf_109_clk _00668_ VGND VGND VPWR VPWR data_array.data0\[7\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10811_ net2428 net984 net507 VGND VGND VPWR VPWR _02556_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11791_ clknet_leaf_237_clk _00599_ VGND VGND VPWR VPWR data_array.data0\[8\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_0_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13530_ clknet_leaf_220_clk _02159_ VGND VGND VPWR VPWR data_array.data1\[0\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_10742_ net1004 net3426 net491 VGND VGND VPWR VPWR _02487_ sky130_fd_sc_hd__mux2_1
XFILLER_13_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10673_ net3030 net1025 net482 VGND VGND VPWR VPWR _02418_ sky130_fd_sc_hd__mux2_1
X_13461_ clknet_leaf_109_clk _02091_ VGND VGND VPWR VPWR tag_array.tag0\[1\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_11_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_173_Right_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12412_ clknet_leaf_70_clk _01106_ VGND VGND VPWR VPWR data_array.data0\[14\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_97_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13392_ clknet_leaf_85_clk _02022_ VGND VGND VPWR VPWR data_array.data1\[8\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12343_ clknet_leaf_267_clk _00017_ VGND VGND VPWR VPWR data_array.rdata0\[25\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_58_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12274_ clknet_leaf_195_clk _01032_ VGND VGND VPWR VPWR tag_array.tag1\[13\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_75_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14013_ clknet_leaf_3_clk _02642_ VGND VGND VPWR VPWR data_array.data1\[5\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
X_11225_ net874 net4416 net655 VGND VGND VPWR VPWR _02968_ sky130_fd_sc_hd__mux2_1
XFILLER_49_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11156_ net893 net4281 net542 VGND VGND VPWR VPWR _02899_ sky130_fd_sc_hd__mux2_1
X_10107_ net2086 net695 net638 VGND VGND VPWR VPWR _01856_ sky130_fd_sc_hd__mux2_1
XFILLER_0_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11087_ net2317 net912 net333 VGND VGND VPWR VPWR _02830_ sky130_fd_sc_hd__mux2_1
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10038_ net934 net2352 net563 VGND VGND VPWR VPWR _01787_ sky130_fd_sc_hd__mux2_1
XFILLER_76_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_762 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_698 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11989_ clknet_leaf_225_clk _00797_ VGND VGND VPWR VPWR data_array.data0\[4\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
X_13728_ clknet_leaf_91_clk _02357_ VGND VGND VPWR VPWR data_array.data1\[1\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_3328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13659_ clknet_leaf_67_clk _02288_ VGND VGND VPWR VPWR data_array.data1\[15\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_83_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06200_ tag_array.tag0\[5\]\[1\] net1593 net1497 tag_array.tag0\[6\]\[1\] VGND VGND
+ VPWR VPWR _03554_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_140_Right_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_171_3653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07180_ data_array.data0\[4\]\[40\] net1412 net1318 data_array.data0\[7\]\[40\] _04444_
+ VGND VGND VPWR VPWR _04445_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_30_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06131_ data_array.rdata0\[46\] net1134 net1113 data_array.rdata1\[46\] VGND VGND
+ VPWR VPWR net303 sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_132_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06062_ fsm.tag_out0\[13\] net1121 _03494_ VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__a21o_1
XFILLER_144_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout406 net408 VGND VGND VPWR VPWR net406 sky130_fd_sc_hd__clkbuf_8
X_09821_ net926 net3517 net386 VGND VGND VPWR VPWR _01572_ sky130_fd_sc_hd__mux2_1
Xfanout417 _05611_ VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__clkbuf_8
XFILLER_141_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout428 net429 VGND VGND VPWR VPWR net428 sky130_fd_sc_hd__buf_4
XFILLER_101_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout439 net441 VGND VGND VPWR VPWR net439 sky130_fd_sc_hd__buf_4
XFILLER_141_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_129_Left_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09752_ net2246 net778 net665 VGND VGND VPWR VPWR _01504_ sky130_fd_sc_hd__mux2_1
X_06964_ data_array.data0\[0\]\[20\] net1412 net1318 data_array.data0\[3\]\[20\] _04248_
+ VGND VGND VPWR VPWR _04249_ sky130_fd_sc_hd__a221o_1
XFILLER_39_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08703_ net3286 net710 net480 VGND VGND VPWR VPWR _00462_ sky130_fd_sc_hd__mux2_1
X_05915_ data_array.rdata0\[28\] net847 net1143 VGND VGND VPWR VPWR _03404_ sky130_fd_sc_hd__o21a_1
X_06895_ data_array.data0\[13\]\[14\] net1570 net1474 data_array.data0\[14\]\[14\]
+ VGND VGND VPWR VPWR _04186_ sky130_fd_sc_hd__a22o_1
X_09683_ net754 net4537 net607 VGND VGND VPWR VPWR _01435_ sky130_fd_sc_hd__mux2_1
X_05846_ data_array.rdata0\[5\] net849 net1144 VGND VGND VPWR VPWR _03358_ sky130_fd_sc_hd__o21a_1
X_08634_ net2144 net787 net511 VGND VGND VPWR VPWR _00393_ sky130_fd_sc_hd__mux2_1
XFILLER_82_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08565_ net695 net4539 net583 VGND VGND VPWR VPWR _00333_ sky130_fd_sc_hd__mux2_1
X_05777_ _03288_ _03290_ _03293_ VGND VGND VPWR VPWR _03294_ sky130_fd_sc_hd__or3_1
X_07516_ net1213 _04745_ _04749_ net1165 VGND VGND VPWR VPWR _04751_ sky130_fd_sc_hd__a22o_1
X_08496_ net1706 net623 VGND VGND VPWR VPWR _00294_ sky130_fd_sc_hd__nand2b_1
XPHY_EDGE_ROW_138_Left_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07447_ data_array.data1\[5\]\[0\] net1556 net1460 data_array.data1\[6\]\[0\] VGND
+ VGND VPWR VPWR _04688_ sky130_fd_sc_hd__a22o_1
XFILLER_167_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_940 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_170_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_170_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_10_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07378_ data_array.data0\[4\]\[58\] net1354 net1260 data_array.data0\[7\]\[58\] _04624_
+ VGND VGND VPWR VPWR _04625_ sky130_fd_sc_hd__a221o_1
XFILLER_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06329_ _03670_ _03671_ VGND VGND VPWR VPWR _00134_ sky130_fd_sc_hd__or2_1
X_09117_ net1074 net4224 net574 VGND VGND VPWR VPWR _00871_ sky130_fd_sc_hd__mux2_1
XFILLER_135_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09048_ net1092 net3328 net415 VGND VGND VPWR VPWR _00802_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_92_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold460 data_array.data1\[2\]\[26\] VGND VGND VPWR VPWR net2111 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_53_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold471 data_array.data0\[10\]\[62\] VGND VGND VPWR VPWR net2122 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_147_Left_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11010_ net2234 net961 net338 VGND VGND VPWR VPWR _02754_ sky130_fd_sc_hd__mux2_1
Xhold482 data_array.data0\[1\]\[61\] VGND VGND VPWR VPWR net2133 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold493 tag_array.tag1\[4\]\[1\] VGND VGND VPWR VPWR net2144 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout940 net941 VGND VGND VPWR VPWR net940 sky130_fd_sc_hd__clkbuf_2
Xfanout951 _05500_ VGND VGND VPWR VPWR net951 sky130_fd_sc_hd__buf_1
Xfanout962 net963 VGND VGND VPWR VPWR net962 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout973 _05488_ VGND VGND VPWR VPWR net973 sky130_fd_sc_hd__buf_1
Xfanout984 _05482_ VGND VGND VPWR VPWR net984 sky130_fd_sc_hd__clkbuf_2
Xfanout995 _05478_ VGND VGND VPWR VPWR net995 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12961_ clknet_leaf_164_clk _01655_ VGND VGND VPWR VPWR tag_array.tag0\[4\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_5_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1160 data_array.data1\[2\]\[52\] VGND VGND VPWR VPWR net2811 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1171 tag_array.tag0\[12\]\[1\] VGND VGND VPWR VPWR net2822 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11912_ clknet_leaf_241_clk _00720_ VGND VGND VPWR VPWR data_array.data0\[5\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1182 tag_array.tag0\[10\]\[2\] VGND VGND VPWR VPWR net2833 sky130_fd_sc_hd__dlygate4sd3_1
X_12892_ clknet_leaf_115_clk _01586_ VGND VGND VPWR VPWR data_array.data0\[12\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1193 data_array.data1\[8\]\[56\] VGND VGND VPWR VPWR net2844 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_16_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ clknet_leaf_20_clk _00651_ VGND VGND VPWR VPWR data_array.data0\[7\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_61_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_68_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_156_Left_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11774_ clknet_leaf_125_clk _00582_ VGND VGND VPWR VPWR data_array.data0\[8\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
X_13513_ clknet_leaf_116_clk _02142_ VGND VGND VPWR VPWR data_array.data1\[0\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_10725_ net1074 net2188 net497 VGND VGND VPWR VPWR _02470_ sky130_fd_sc_hd__mux2_1
XFILLER_41_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_161_clk clknet_5_25__leaf_clk VGND VGND VPWR VPWR clknet_leaf_161_clk
+ sky130_fd_sc_hd__clkbuf_8
X_14493_ clknet_leaf_161_clk _03116_ VGND VGND VPWR VPWR tag_array.dirty0\[12\] sky130_fd_sc_hd__dfxtp_1
X_13444_ clknet_leaf_105_clk _02074_ VGND VGND VPWR VPWR tag_array.tag0\[1\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_10656_ net2218 net1094 net484 VGND VGND VPWR VPWR _02401_ sky130_fd_sc_hd__mux2_1
XFILLER_16_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload16 clknet_leaf_1_clk VGND VGND VPWR VPWR clkload16/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_70_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload27 clknet_leaf_266_clk VGND VGND VPWR VPWR clkload27/Y sky130_fd_sc_hd__clkinv_8
X_10587_ net858 net2652 net457 VGND VGND VPWR VPWR _02332_ sky130_fd_sc_hd__mux2_1
X_13375_ clknet_leaf_168_clk _02005_ VGND VGND VPWR VPWR tag_array.tag0\[2\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload38 clknet_leaf_8_clk VGND VGND VPWR VPWR clkload38/Y sky130_fd_sc_hd__clkinv_2
XFILLER_103_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload49 clknet_leaf_259_clk VGND VGND VPWR VPWR clkload49/Y sky130_fd_sc_hd__bufinv_16
XFILLER_86_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12326_ clknet_leaf_15_clk _00062_ VGND VGND VPWR VPWR data_array.rdata0\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_55_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_165_Left_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12257_ clknet_leaf_231_clk _01015_ VGND VGND VPWR VPWR tag_array.tag1\[14\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_107_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11208_ net943 net4409 net657 VGND VGND VPWR VPWR _02951_ sky130_fd_sc_hd__mux2_1
X_12188_ clknet_leaf_171_clk _00996_ VGND VGND VPWR VPWR tag_array.tag0\[14\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_96_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_147_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11139_ net960 net2390 net545 VGND VGND VPWR VPWR _02882_ sky130_fd_sc_hd__mux2_1
XFILLER_1_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_147_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_802 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_1044 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05700_ _03214_ _03215_ _03216_ VGND VGND VPWR VPWR _03217_ sky130_fd_sc_hd__or3_1
XFILLER_23_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06680_ net1181 _03985_ _03989_ net1229 VGND VGND VPWR VPWR _03991_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_125_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05631_ fsm.lru_out fsm.valid1 dirty_way1 _03149_ VGND VGND VPWR VPWR _03150_ sky130_fd_sc_hd__a31o_1
XFILLER_93_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08350_ net1123 _05469_ VGND VGND VPWR VPWR _05470_ sky130_fd_sc_hd__and2_1
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07301_ data_array.data0\[4\]\[51\] net1332 net1238 data_array.data0\[7\]\[51\] _04554_
+ VGND VGND VPWR VPWR _04555_ sky130_fd_sc_hd__a221o_1
XFILLER_149_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08281_ net1125 _05423_ VGND VGND VPWR VPWR _05424_ sky130_fd_sc_hd__and2_1
XFILLER_60_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_152_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_152_clk
+ sky130_fd_sc_hd__clkbuf_8
X_07232_ data_array.data0\[13\]\[45\] net1535 net1439 data_array.data0\[14\]\[45\]
+ VGND VGND VPWR VPWR _04492_ sky130_fd_sc_hd__a22o_1
XFILLER_118_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07163_ net1631 _04423_ _04427_ net1205 VGND VGND VPWR VPWR _04430_ sky130_fd_sc_hd__a22o_1
XFILLER_9_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06114_ data_array.rdata0\[29\] net1140 net1114 data_array.rdata1\[29\] VGND VGND
+ VPWR VPWR net284 sky130_fd_sc_hd__a22o_1
XFILLER_161_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07094_ data_array.data0\[8\]\[32\] net1333 net1239 data_array.data0\[11\]\[32\]
+ _04366_ VGND VGND VPWR VPWR _04367_ sky130_fd_sc_hd__a221o_1
XFILLER_105_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06045_ net1163 net4 fsm.tag_out1\[5\] net1132 VGND VGND VPWR VPWR _03486_ sky130_fd_sc_hd__a22o_1
XFILLER_120_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_184_3888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09804_ net993 net2973 net391 VGND VGND VPWR VPWR _01555_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_184_3899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07996_ data_array.data1\[12\]\[50\] net1337 net1243 data_array.data1\[15\]\[50\]
+ _05186_ VGND VGND VPWR VPWR _05187_ sky130_fd_sc_hd__a221o_1
XFILLER_74_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09735_ net747 net2713 net680 VGND VGND VPWR VPWR _01487_ sky130_fd_sc_hd__mux2_1
X_06947_ data_array.data0\[12\]\[19\] net1390 net1296 data_array.data0\[15\]\[19\]
+ _04232_ VGND VGND VPWR VPWR _04233_ sky130_fd_sc_hd__a221o_1
XFILLER_74_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09666_ net722 net3588 net613 VGND VGND VPWR VPWR _01418_ sky130_fd_sc_hd__mux2_1
X_06878_ net1225 _04165_ _04169_ net1177 VGND VGND VPWR VPWR _04171_ sky130_fd_sc_hd__a22o_1
XFILLER_28_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08617_ net756 net4622 net523 VGND VGND VPWR VPWR _00376_ sky130_fd_sc_hd__mux2_1
XFILLER_15_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05829_ _03309_ _03343_ _03344_ _03345_ VGND VGND VPWR VPWR _03346_ sky130_fd_sc_hd__or4_1
X_09597_ net961 net3789 net396 VGND VGND VPWR VPWR _01349_ sky130_fd_sc_hd__mux2_1
XFILLER_27_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08548_ net765 net3733 net588 VGND VGND VPWR VPWR _00316_ sky130_fd_sc_hd__mux2_1
XFILLER_70_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08479_ _03507_ _03514_ VGND VGND VPWR VPWR _05556_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_143_clk clknet_5_30__leaf_clk VGND VGND VPWR VPWR clknet_leaf_143_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_11_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10510_ net905 net3646 net344 VGND VGND VPWR VPWR _02255_ sky130_fd_sc_hd__mux2_1
X_11490_ clknet_leaf_155_clk _00299_ VGND VGND VPWR VPWR tag_array.valid0\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_168_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10441_ net1904 net890 net663 VGND VGND VPWR VPWR _02187_ sky130_fd_sc_hd__mux2_1
XFILLER_148_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13160_ clknet_leaf_196_clk _01854_ VGND VGND VPWR VPWR tag_array.tag1\[8\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_10372_ net713 net2249 net538 VGND VGND VPWR VPWR _02119_ sky130_fd_sc_hd__mux2_1
XFILLER_108_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12111_ clknet_leaf_239_clk _00919_ VGND VGND VPWR VPWR data_array.data1\[14\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
X_13091_ clknet_leaf_84_clk _01785_ VGND VGND VPWR VPWR data_array.data1\[13\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_152_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12042_ clknet_leaf_208_clk _00850_ VGND VGND VPWR VPWR data_array.data0\[6\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_123_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold290 tag_array.tag1\[0\]\[8\] VGND VGND VPWR VPWR net1941 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout770 net771 VGND VGND VPWR VPWR net770 sky130_fd_sc_hd__clkbuf_2
Xfanout781 _05371_ VGND VGND VPWR VPWR net781 sky130_fd_sc_hd__clkbuf_2
XFILLER_172_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout792 _05365_ VGND VGND VPWR VPWR net792 sky130_fd_sc_hd__buf_1
X_13993_ clknet_leaf_74_clk _02622_ VGND VGND VPWR VPWR data_array.data1\[5\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
X_12944_ clknet_leaf_57_clk _01638_ VGND VGND VPWR VPWR data_array.data0\[13\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_142_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12875_ clknet_leaf_47_clk _01569_ VGND VGND VPWR VPWR data_array.data0\[12\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_73_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ clknet_leaf_30_clk _00634_ VGND VGND VPWR VPWR data_array.data0\[7\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_83_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_134_clk clknet_5_31__leaf_clk VGND VGND VPWR VPWR clknet_leaf_134_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11757_ clknet_leaf_191_clk _00565_ VGND VGND VPWR VPWR data_array.data0\[8\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_10708_ net2571 net886 net479 VGND VGND VPWR VPWR _02453_ sky130_fd_sc_hd__mux2_1
XFILLER_119_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14476_ clknet_leaf_120_clk _03099_ VGND VGND VPWR VPWR data_array.data1\[7\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_147_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11688_ clknet_leaf_194_clk _00496_ VGND VGND VPWR VPWR tag_array.tag1\[15\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_174_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13427_ clknet_leaf_79_clk _02057_ VGND VGND VPWR VPWR data_array.data1\[8\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload105 clknet_leaf_90_clk VGND VGND VPWR VPWR clkload105/Y sky130_fd_sc_hd__inv_8
X_10639_ net2027 net906 net466 VGND VGND VPWR VPWR _02384_ sky130_fd_sc_hd__mux2_1
Xclkload116 clknet_leaf_72_clk VGND VGND VPWR VPWR clkload116/Y sky130_fd_sc_hd__inv_6
Xclkload127 clknet_leaf_82_clk VGND VGND VPWR VPWR clkload127/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_10_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload138 clknet_leaf_220_clk VGND VGND VPWR VPWR clkload138/Y sky130_fd_sc_hd__inv_8
Xclkload149 clknet_leaf_167_clk VGND VGND VPWR VPWR clkload149/Y sky130_fd_sc_hd__clkinv_4
XFILLER_6_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13358_ clknet_leaf_176_clk _01988_ VGND VGND VPWR VPWR tag_array.tag0\[2\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_114_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12309_ clknet_leaf_136_clk _01067_ VGND VGND VPWR VPWR tag_array.tag1\[12\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_149_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13289_ clknet_leaf_124_clk _01919_ VGND VGND VPWR VPWR data_array.data0\[11\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_149_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_3552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2608 tag_array.tag0\[15\]\[6\] VGND VGND VPWR VPWR net4259 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2619 tag_array.tag1\[13\]\[7\] VGND VGND VPWR VPWR net4270 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_68_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07850_ data_array.data1\[1\]\[37\] net1544 net1448 data_array.data1\[2\]\[37\] VGND
+ VGND VPWR VPWR _05054_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_127_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1907 tag_array.tag1\[13\]\[13\] VGND VGND VPWR VPWR net3558 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_127_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1918 data_array.data0\[9\]\[37\] VGND VGND VPWR VPWR net3569 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06801_ net1219 _04095_ _04099_ net1171 VGND VGND VPWR VPWR _04101_ sky130_fd_sc_hd__a22o_1
Xhold1929 data_array.data0\[11\]\[18\] VGND VGND VPWR VPWR net3580 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07781_ _04990_ _04991_ VGND VGND VPWR VPWR _00087_ sky130_fd_sc_hd__or2_1
Xinput3 cpu_addr[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_2
X_09520_ net748 net3676 net622 VGND VGND VPWR VPWR _01273_ sky130_fd_sc_hd__mux2_1
X_06732_ tag_array.tag1\[1\]\[24\] net1562 net1466 tag_array.tag1\[2\]\[24\] VGND
+ VGND VPWR VPWR _04038_ sky130_fd_sc_hd__a22o_1
XFILLER_37_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09451_ net863 net2654 net588 VGND VGND VPWR VPWR _01204_ sky130_fd_sc_hd__mux2_1
X_06663_ tag_array.tag1\[0\]\[18\] net1372 net1278 tag_array.tag1\[3\]\[18\] _03974_
+ VGND VGND VPWR VPWR _03975_ sky130_fd_sc_hd__a221o_1
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05614_ net32 VGND VGND VPWR VPWR _03136_ sky130_fd_sc_hd__inv_2
X_08402_ net2034 net941 net693 VGND VGND VPWR VPWR _00263_ sky130_fd_sc_hd__mux2_1
X_06594_ tag_array.tag1\[13\]\[12\] net1558 net1462 tag_array.tag1\[14\]\[12\] VGND
+ VGND VPWR VPWR _03912_ sky130_fd_sc_hd__a22o_1
X_09382_ net872 net4443 net406 VGND VGND VPWR VPWR _01135_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08333_ net1933 net1033 net691 VGND VGND VPWR VPWR _00240_ sky130_fd_sc_hd__mux2_1
XFILLER_51_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_125_clk clknet_5_27__leaf_clk VGND VGND VPWR VPWR clknet_leaf_125_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_178_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08264_ fsm.tag_out1\[23\] net817 net809 fsm.tag_out0\[23\] _05410_ VGND VGND VPWR
+ VPWR _05411_ sky130_fd_sc_hd__a221o_2
XFILLER_20_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07215_ data_array.data0\[12\]\[43\] net1377 net1283 data_array.data0\[15\]\[43\]
+ _04476_ VGND VGND VPWR VPWR _04477_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_41_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08195_ fsm.tag_out1\[0\] net817 net809 fsm.tag_out0\[0\] _05363_ VGND VGND VPWR
+ VPWR _05365_ sky130_fd_sc_hd__a221o_4
XTAP_TAPCELL_ROW_41_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07146_ data_array.data0\[1\]\[37\] net1546 net1450 data_array.data0\[2\]\[37\] VGND
+ VGND VPWR VPWR _04414_ sky130_fd_sc_hd__a22o_1
XFILLER_106_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07077_ _04350_ _04351_ VGND VGND VPWR VPWR _00023_ sky130_fd_sc_hd__or2_1
XFILLER_156_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06028_ _03476_ net1137 VGND VGND VPWR VPWR _03478_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_7_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1009 net1010 VGND VGND VPWR VPWR net1009 sky130_fd_sc_hd__clkbuf_2
XFILLER_99_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07979_ _05170_ _05171_ VGND VGND VPWR VPWR _00106_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_87_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_87_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09718_ net716 net3656 net610 VGND VGND VPWR VPWR _01470_ sky130_fd_sc_hd__mux2_1
X_10990_ net2057 net1042 net339 VGND VGND VPWR VPWR _02734_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09649_ net793 net2875 net613 VGND VGND VPWR VPWR _01401_ sky130_fd_sc_hd__mux2_1
XFILLER_15_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12660_ clknet_leaf_87_clk _01354_ VGND VGND VPWR VPWR data_array.data0\[15\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ clknet_leaf_233_clk _00419_ VGND VGND VPWR VPWR tag_array.tag1\[3\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_26_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_116_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_116_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12591_ clknet_leaf_142_clk _01285_ VGND VGND VPWR VPWR tag_array.tag0\[10\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14330_ clknet_leaf_242_clk _02959_ VGND VGND VPWR VPWR data_array.data1\[11\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_61_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11542_ clknet_leaf_141_clk _00350_ VGND VGND VPWR VPWR tag_array.tag1\[6\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14261_ clknet_leaf_28_clk _02890_ VGND VGND VPWR VPWR data_array.data1\[12\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
X_11473_ clknet_leaf_110_clk _00283_ VGND VGND VPWR VPWR data_array.data0\[0\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13212_ clknet_leaf_53_clk _00107_ VGND VGND VPWR VPWR data_array.rdata1\[49\] sky130_fd_sc_hd__dfxtp_1
X_10424_ net2100 net958 net669 VGND VGND VPWR VPWR _02170_ sky130_fd_sc_hd__mux2_1
XFILLER_171_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14192_ clknet_leaf_109_clk _02821_ VGND VGND VPWR VPWR data_array.data0\[2\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13143_ clknet_leaf_134_clk _01837_ VGND VGND VPWR VPWR tag_array.tag1\[8\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_10355_ _05371_ net3610 net538 VGND VGND VPWR VPWR _02102_ sky130_fd_sc_hd__mux2_1
X_10286_ net3357 net1017 net637 VGND VGND VPWR VPWR _02033_ sky130_fd_sc_hd__mux2_1
X_13074_ clknet_leaf_263_clk _01768_ VGND VGND VPWR VPWR data_array.data1\[13\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_112_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1510 net1516 VGND VGND VPWR VPWR net1510 sky130_fd_sc_hd__buf_2
X_12025_ clknet_leaf_243_clk _00833_ VGND VGND VPWR VPWR data_array.data0\[6\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout1521 net1543 VGND VGND VPWR VPWR net1521 sky130_fd_sc_hd__clkbuf_2
Xfanout1532 net1533 VGND VGND VPWR VPWR net1532 sky130_fd_sc_hd__clkbuf_4
Xfanout1543 _03508_ VGND VGND VPWR VPWR net1543 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_144_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1554 net1566 VGND VGND VPWR VPWR net1554 sky130_fd_sc_hd__buf_2
XFILLER_120_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1565 net1566 VGND VGND VPWR VPWR net1565 sky130_fd_sc_hd__buf_2
Xfanout1576 net1591 VGND VGND VPWR VPWR net1576 sky130_fd_sc_hd__clkbuf_4
Xfanout1587 net1591 VGND VGND VPWR VPWR net1587 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_161_3460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1598 net1599 VGND VGND VPWR VPWR net1598 sky130_fd_sc_hd__clkbuf_4
X_13976_ clknet_leaf_214_clk _02605_ VGND VGND VPWR VPWR data_array.data1\[5\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_122_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12927_ clknet_leaf_97_clk _01621_ VGND VGND VPWR VPWR data_array.data0\[13\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12858_ clknet_leaf_247_clk _01552_ VGND VGND VPWR VPWR data_array.data0\[12\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_476 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11809_ clknet_leaf_45_clk _00617_ VGND VGND VPWR VPWR data_array.data0\[7\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_107_clk clknet_5_25__leaf_clk VGND VGND VPWR VPWR clknet_leaf_107_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12789_ clknet_leaf_133_clk _01483_ VGND VGND VPWR VPWR tag_array.tag1\[10\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14459_ clknet_leaf_45_clk _03082_ VGND VGND VPWR VPWR data_array.data1\[7\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
X_07000_ _04280_ _04281_ VGND VGND VPWR VPWR _00015_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08951_ net961 net3741 net428 VGND VGND VPWR VPWR _00707_ sky130_fd_sc_hd__mux2_1
XFILLER_103_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2405 tag_array.tag1\[5\]\[3\] VGND VGND VPWR VPWR net4056 sky130_fd_sc_hd__dlygate4sd3_1
X_07902_ _05100_ _05101_ VGND VGND VPWR VPWR _00099_ sky130_fd_sc_hd__or2_1
Xhold2416 data_array.data1\[12\]\[18\] VGND VGND VPWR VPWR net4067 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2427 data_array.data1\[9\]\[38\] VGND VGND VPWR VPWR net4078 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_181_3836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08882_ net976 net2520 net438 VGND VGND VPWR VPWR _00639_ sky130_fd_sc_hd__mux2_1
Xhold2438 data_array.data1\[7\]\[36\] VGND VGND VPWR VPWR net4089 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1704 data_array.data1\[5\]\[27\] VGND VGND VPWR VPWR net3355 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2449 tag_array.tag0\[1\]\[14\] VGND VGND VPWR VPWR net4100 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_102_Left_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1715 tag_array.tag0\[15\]\[24\] VGND VGND VPWR VPWR net3366 sky130_fd_sc_hd__dlygate4sd3_1
X_07833_ data_array.data1\[0\]\[35\] net1335 net1241 data_array.data1\[3\]\[35\] _05038_
+ VGND VGND VPWR VPWR _05039_ sky130_fd_sc_hd__a221o_1
XFILLER_57_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1726 tag_array.tag0\[2\]\[20\] VGND VGND VPWR VPWR net3377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1737 tag_array.tag1\[15\]\[23\] VGND VGND VPWR VPWR net3388 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1748 data_array.data1\[13\]\[24\] VGND VGND VPWR VPWR net3399 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_81_Right_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_5_25__f_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_5_25__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_38_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1759 data_array.data0\[6\]\[12\] VGND VGND VPWR VPWR net3410 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_568 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07764_ data_array.data1\[9\]\[29\] net1578 net1482 data_array.data1\[10\]\[29\]
+ VGND VGND VPWR VPWR _04976_ sky130_fd_sc_hd__a22o_1
XFILLER_72_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09503_ net716 net4540 net625 VGND VGND VPWR VPWR _01256_ sky130_fd_sc_hd__mux2_1
X_06715_ tag_array.tag1\[9\]\[23\] net1610 net1514 tag_array.tag1\[10\]\[23\] VGND
+ VGND VPWR VPWR _04022_ sky130_fd_sc_hd__a22o_1
XFILLER_25_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07695_ data_array.data1\[12\]\[23\] net1359 net1265 data_array.data1\[15\]\[23\]
+ _04912_ VGND VGND VPWR VPWR _04913_ sky130_fd_sc_hd__a221o_1
X_09434_ net931 net2342 net580 VGND VGND VPWR VPWR _01187_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_179_3798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06646_ net1210 _03953_ _03957_ net1636 VGND VGND VPWR VPWR _03960_ sky130_fd_sc_hd__a22o_1
XFILLER_25_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09365_ net941 net4523 net409 VGND VGND VPWR VPWR _01118_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06577_ tag_array.tag1\[8\]\[10\] net1404 net1310 tag_array.tag1\[11\]\[10\] _03896_
+ VGND VGND VPWR VPWR _03897_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_111_Left_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08316_ net104 net39 net1640 VGND VGND VPWR VPWR _05447_ sky130_fd_sc_hd__mux2_1
X_09296_ net695 net2807 net559 VGND VGND VPWR VPWR _01050_ sky130_fd_sc_hd__mux2_1
XANTENNA_30 _05551_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_41 net508 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_52 net1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_90_Right_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_63 net1543 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08247_ net724 net4010 net804 VGND VGND VPWR VPWR _00213_ sky130_fd_sc_hd__mux2_1
XANTENNA_74 _03480_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_85 net1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_506 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08178_ net4614 net849 _03285_ VGND VGND VPWR VPWR _00185_ sky130_fd_sc_hd__and3_1
XFILLER_21_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07129_ data_array.data0\[0\]\[35\] net1337 net1243 data_array.data0\[3\]\[35\] _04398_
+ VGND VGND VPWR VPWR _04399_ sky130_fd_sc_hd__a221o_1
XFILLER_122_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10140_ net986 net4274 net366 VGND VGND VPWR VPWR _01888_ sky130_fd_sc_hd__mux2_1
XFILLER_0_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput170 net170 VGND VGND VPWR VPWR cpu_rdata[14] sky130_fd_sc_hd__buf_6
Xoutput181 net181 VGND VGND VPWR VPWR cpu_rdata[24] sky130_fd_sc_hd__buf_6
XFILLER_0_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput192 net192 VGND VGND VPWR VPWR cpu_rdata[34] sky130_fd_sc_hd__buf_2
X_10071_ net739 net3099 net601 VGND VGND VPWR VPWR _01820_ sky130_fd_sc_hd__mux2_1
XFILLER_88_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2950 data_array.data0\[9\]\[1\] VGND VGND VPWR VPWR net4601 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2961 data_array.data1\[3\]\[33\] VGND VGND VPWR VPWR net4612 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2972 data_array.data1\[11\]\[23\] VGND VGND VPWR VPWR net4623 sky130_fd_sc_hd__dlygate4sd3_1
X_13830_ clknet_leaf_120_clk _02459_ VGND VGND VPWR VPWR data_array.data1\[2\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13761_ clknet_leaf_249_clk _02390_ VGND VGND VPWR VPWR data_array.data1\[1\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
X_10973_ net2606 net1108 net340 VGND VGND VPWR VPWR _02717_ sky130_fd_sc_hd__mux2_1
XFILLER_44_966 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12712_ clknet_leaf_143_clk _01406_ VGND VGND VPWR VPWR tag_array.tag0\[7\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_100_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13692_ clknet_leaf_208_clk _02321_ VGND VGND VPWR VPWR data_array.data1\[15\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12643_ clknet_leaf_262_clk _01337_ VGND VGND VPWR VPWR data_array.data0\[15\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_80_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12574_ clknet_leaf_179_clk _01268_ VGND VGND VPWR VPWR tag_array.tag0\[10\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_129_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_885 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14313_ clknet_leaf_77_clk _02942_ VGND VGND VPWR VPWR data_array.data1\[11\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
X_11525_ clknet_leaf_188_clk _00333_ VGND VGND VPWR VPWR tag_array.tag1\[9\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14244_ clknet_leaf_30_clk _02873_ VGND VGND VPWR VPWR data_array.data1\[12\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11456_ clknet_leaf_20_clk _00266_ VGND VGND VPWR VPWR data_array.data0\[0\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_78_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10407_ net2372 net1025 net665 VGND VGND VPWR VPWR _02153_ sky130_fd_sc_hd__mux2_1
X_14175_ clknet_leaf_225_clk _02804_ VGND VGND VPWR VPWR data_array.data0\[2\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_78_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11387_ clknet_leaf_167_clk _00197_ VGND VGND VPWR VPWR tag_array.tag1\[7\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13126_ clknet_leaf_139_clk _01820_ VGND VGND VPWR VPWR tag_array.tag0\[3\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_180_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10338_ net748 net3587 net592 VGND VGND VPWR VPWR _02085_ sky130_fd_sc_hd__mux2_1
XFILLER_140_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_163_3500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13057_ clknet_leaf_19_clk _01751_ VGND VGND VPWR VPWR data_array.data1\[13\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_111_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10269_ net2824 net1087 net633 VGND VGND VPWR VPWR _02016_ sky130_fd_sc_hd__mux2_1
Xfanout1340 net1342 VGND VGND VPWR VPWR net1340 sky130_fd_sc_hd__clkbuf_4
X_12008_ clknet_leaf_15_clk _00816_ VGND VGND VPWR VPWR data_array.data0\[6\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout1351 net1352 VGND VGND VPWR VPWR net1351 sky130_fd_sc_hd__clkbuf_2
Xfanout1362 net1363 VGND VGND VPWR VPWR net1362 sky130_fd_sc_hd__clkbuf_4
Xfanout1373 net1375 VGND VGND VPWR VPWR net1373 sky130_fd_sc_hd__clkbuf_4
XFILLER_66_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1384 net1385 VGND VGND VPWR VPWR net1384 sky130_fd_sc_hd__clkbuf_4
Xfanout1395 net1399 VGND VGND VPWR VPWR net1395 sky130_fd_sc_hd__clkbuf_4
XFILLER_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13959_ clknet_leaf_204_clk _02588_ VGND VGND VPWR VPWR data_array.data1\[4\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06500_ tag_array.tag1\[12\]\[3\] net1371 net1277 tag_array.tag1\[15\]\[3\] _03826_
+ VGND VGND VPWR VPWR _03827_ sky130_fd_sc_hd__a221o_1
X_07480_ data_array.data1\[1\]\[3\] net1574 net1478 data_array.data1\[2\]\[3\] VGND
+ VGND VPWR VPWR _04718_ sky130_fd_sc_hd__a22o_1
XFILLER_50_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06431_ tag_array.tag0\[5\]\[22\] net1565 net1469 tag_array.tag0\[6\]\[22\] VGND
+ VGND VPWR VPWR _03764_ sky130_fd_sc_hd__a22o_1
X_09150_ net943 net4084 net575 VGND VGND VPWR VPWR _00904_ sky130_fd_sc_hd__mux2_1
XFILLER_148_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06362_ _03700_ _03701_ VGND VGND VPWR VPWR _00137_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_174_3695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08101_ data_array.data1\[9\]\[60\] net1604 net1508 data_array.data1\[10\]\[60\]
+ VGND VGND VPWR VPWR _05282_ sky130_fd_sc_hd__a22o_1
X_09081_ net961 net2907 net412 VGND VGND VPWR VPWR _00835_ sky130_fd_sc_hd__mux2_1
X_06293_ tag_array.tag0\[4\]\[9\] net1409 net1315 tag_array.tag0\[7\]\[9\] _03638_
+ VGND VGND VPWR VPWR _03639_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_135_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08032_ net1615 _05213_ _05217_ net1189 VGND VGND VPWR VPWR _05220_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_135_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput50 cpu_wdata[24] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_1
Xinput61 cpu_wdata[34] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_1
Xinput72 cpu_wdata[44] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_1
Xhold801 data_array.data0\[4\]\[28\] VGND VGND VPWR VPWR net2452 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_174_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold812 tag_array.tag1\[4\]\[22\] VGND VGND VPWR VPWR net2463 sky130_fd_sc_hd__dlygate4sd3_1
Xinput83 cpu_wdata[54] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_1
Xhold823 data_array.data1\[10\]\[9\] VGND VGND VPWR VPWR net2474 sky130_fd_sc_hd__dlygate4sd3_1
Xinput94 cpu_wdata[6] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_1
Xhold834 data_array.data0\[14\]\[31\] VGND VGND VPWR VPWR net2485 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold845 data_array.data0\[0\]\[63\] VGND VGND VPWR VPWR net2496 sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 data_array.data1\[15\]\[31\] VGND VGND VPWR VPWR net2507 sky130_fd_sc_hd__dlygate4sd3_1
Xhold867 data_array.data0\[6\]\[15\] VGND VGND VPWR VPWR net2518 sky130_fd_sc_hd__dlygate4sd3_1
Xhold878 data_array.data1\[10\]\[14\] VGND VGND VPWR VPWR net2529 sky130_fd_sc_hd__dlygate4sd3_1
Xhold889 data_array.data1\[11\]\[62\] VGND VGND VPWR VPWR net2540 sky130_fd_sc_hd__dlygate4sd3_1
X_09983_ net896 net4356 net370 VGND VGND VPWR VPWR _01732_ sky130_fd_sc_hd__mux2_1
Xhold2202 tag_array.tag0\[4\]\[13\] VGND VGND VPWR VPWR net3853 sky130_fd_sc_hd__dlygate4sd3_1
X_08934_ net1028 net4587 net432 VGND VGND VPWR VPWR _00690_ sky130_fd_sc_hd__mux2_1
XFILLER_131_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2213 tag_array.tag0\[1\]\[10\] VGND VGND VPWR VPWR net3864 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2224 data_array.data0\[10\]\[17\] VGND VGND VPWR VPWR net3875 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_36_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2235 tag_array.tag1\[9\]\[11\] VGND VGND VPWR VPWR net3886 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2246 data_array.data1\[9\]\[57\] VGND VGND VPWR VPWR net3897 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1501 tag_array.tag0\[10\]\[3\] VGND VGND VPWR VPWR net3152 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1512 data_array.data1\[12\]\[60\] VGND VGND VPWR VPWR net3163 sky130_fd_sc_hd__dlygate4sd3_1
X_08865_ net1047 net4324 net436 VGND VGND VPWR VPWR _00622_ sky130_fd_sc_hd__mux2_1
Xhold2257 data_array.data0\[3\]\[32\] VGND VGND VPWR VPWR net3908 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1523 data_array.data0\[15\]\[58\] VGND VGND VPWR VPWR net3174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2268 tag_array.tag0\[4\]\[5\] VGND VGND VPWR VPWR net3919 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1534 data_array.data1\[5\]\[4\] VGND VGND VPWR VPWR net3185 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2279 data_array.data1\[1\]\[24\] VGND VGND VPWR VPWR net3930 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1545 data_array.data1\[12\]\[58\] VGND VGND VPWR VPWR net3196 sky130_fd_sc_hd__dlygate4sd3_1
X_07816_ data_array.data1\[12\]\[34\] net1341 net1247 data_array.data1\[15\]\[34\]
+ _05022_ VGND VGND VPWR VPWR _05023_ sky130_fd_sc_hd__a221o_1
Xhold1556 data_array.data0\[8\]\[0\] VGND VGND VPWR VPWR net3207 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_84_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1567 data_array.data0\[10\]\[3\] VGND VGND VPWR VPWR net3218 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08796_ net2131 net1060 net448 VGND VGND VPWR VPWR _00554_ sky130_fd_sc_hd__mux2_1
Xhold1578 tag_array.tag0\[11\]\[21\] VGND VGND VPWR VPWR net3229 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_28_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1589 tag_array.tag1\[1\]\[10\] VGND VGND VPWR VPWR net3240 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_28_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07747_ net1218 _04955_ _04959_ net1170 VGND VGND VPWR VPWR _04961_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_154_Right_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07678_ data_array.data1\[5\]\[21\] net1555 net1459 data_array.data1\[6\]\[21\] VGND
+ VGND VPWR VPWR _04898_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09417_ net998 net4511 net581 VGND VGND VPWR VPWR _01170_ sky130_fd_sc_hd__mux2_1
X_06629_ tag_array.tag1\[1\]\[15\] net1576 net1480 tag_array.tag1\[2\]\[15\] VGND
+ VGND VPWR VPWR _03944_ sky130_fd_sc_hd__a22o_1
XFILLER_13_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09348_ net1010 net3303 net402 VGND VGND VPWR VPWR _01101_ sky130_fd_sc_hd__mux2_1
XFILLER_166_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09279_ net765 net4270 net565 VGND VGND VPWR VPWR _01033_ sky130_fd_sc_hd__mux2_1
X_11310_ net1054 net3476 net800 VGND VGND VPWR VPWR _03053_ sky130_fd_sc_hd__mux2_1
XFILLER_148_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12290_ clknet_leaf_196_clk _01048_ VGND VGND VPWR VPWR tag_array.tag1\[13\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_1013 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11241_ net1066 net3697 net685 VGND VGND VPWR VPWR _02984_ sky130_fd_sc_hd__mux2_1
XFILLER_107_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11172_ net1087 net4482 net648 VGND VGND VPWR VPWR _02915_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10123_ net1053 net4481 net366 VGND VGND VPWR VPWR _01871_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_73_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_971 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10054_ net870 net3015 net564 VGND VGND VPWR VPWR _01803_ sky130_fd_sc_hd__mux2_1
XFILLER_57_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2780 data_array.data0\[14\]\[51\] VGND VGND VPWR VPWR net4431 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_180_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2791 data_array.data1\[15\]\[51\] VGND VGND VPWR VPWR net4442 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13813_ clknet_leaf_26_clk _02442_ VGND VGND VPWR VPWR data_array.data1\[2\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_180_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_121_Right_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13744_ clknet_leaf_123_clk _02373_ VGND VGND VPWR VPWR data_array.data1\[1\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_44_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10956_ net918 net3901 net532 VGND VGND VPWR VPWR _02701_ sky130_fd_sc_hd__mux2_1
XFILLER_32_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_139_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13675_ clknet_leaf_259_clk _02304_ VGND VGND VPWR VPWR data_array.data1\[15\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
X_10887_ net937 net2346 net519 VGND VGND VPWR VPWR _02632_ sky130_fd_sc_hd__mux2_1
XFILLER_31_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12626_ clknet_leaf_18_clk _01320_ VGND VGND VPWR VPWR data_array.data0\[15\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_156_3370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12557_ clknet_leaf_173_clk _01251_ VGND VGND VPWR VPWR tag_array.tag0\[11\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_117_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_152_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11508_ clknet_leaf_134_clk _00316_ VGND VGND VPWR VPWR tag_array.tag1\[9\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_152_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12488_ clknet_leaf_122_clk _01182_ VGND VGND VPWR VPWR data_array.data1\[9\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_176_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold108 tag_array.tag1\[4\]\[16\] VGND VGND VPWR VPWR net1759 sky130_fd_sc_hd__dlygate4sd3_1
Xhold119 data_array.data1\[4\]\[17\] VGND VGND VPWR VPWR net1770 sky130_fd_sc_hd__dlygate4sd3_1
X_14227_ clknet_leaf_35_clk _02856_ VGND VGND VPWR VPWR data_array.data1\[12\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_113_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11439_ clknet_leaf_29_clk _00249_ VGND VGND VPWR VPWR data_array.data0\[0\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_171_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14158_ clknet_leaf_270_clk _02787_ VGND VGND VPWR VPWR data_array.data0\[2\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_130_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13109_ clknet_leaf_119_clk _01803_ VGND VGND VPWR VPWR data_array.data1\[13\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
X_14089_ clknet_leaf_262_clk _02718_ VGND VGND VPWR VPWR data_array.data0\[1\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_06980_ data_array.data0\[8\]\[22\] net1342 net1248 data_array.data0\[11\]\[22\]
+ _04262_ VGND VGND VPWR VPWR _04263_ sky130_fd_sc_hd__a221o_1
XFILLER_140_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05931_ data_array.rdata1\[33\] net832 net841 VGND VGND VPWR VPWR _03415_ sky130_fd_sc_hd__a21o_1
XFILLER_112_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1170 net1174 VGND VGND VPWR VPWR net1170 sky130_fd_sc_hd__buf_4
X_08650_ net2217 net724 net510 VGND VGND VPWR VPWR _00409_ sky130_fd_sc_hd__mux2_1
Xfanout1181 net1182 VGND VGND VPWR VPWR net1181 sky130_fd_sc_hd__clkbuf_4
X_05862_ data_array.rdata1\[10\] net1657 net843 VGND VGND VPWR VPWR _03369_ sky130_fd_sc_hd__a21o_1
Xfanout1192 net1194 VGND VGND VPWR VPWR net1192 sky130_fd_sc_hd__buf_4
X_07601_ data_array.data1\[1\]\[14\] net1567 net1471 data_array.data1\[2\]\[14\] VGND
+ VGND VPWR VPWR _04828_ sky130_fd_sc_hd__a22o_1
XFILLER_26_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08581_ net822 net813 net854 _05590_ VGND VGND VPWR VPWR _05606_ sky130_fd_sc_hd__or4b_4
X_05793_ _03140_ fsm.tag_out1\[14\] _03279_ VGND VGND VPWR VPWR _03310_ sky130_fd_sc_hd__a21o_1
X_07532_ data_array.data1\[4\]\[8\] net1344 net1250 data_array.data1\[7\]\[8\] _04764_
+ VGND VGND VPWR VPWR _04765_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_176_3735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_176_3746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07463_ data_array.data1\[13\]\[2\] net1526 net1430 data_array.data1\[14\]\[2\] VGND
+ VGND VPWR VPWR _04702_ sky130_fd_sc_hd__a22o_1
XFILLER_179_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09202_ net770 net3766 net632 VGND VGND VPWR VPWR _00956_ sky130_fd_sc_hd__mux2_1
XFILLER_22_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06414_ tag_array.tag0\[0\]\[20\] net1368 net1274 tag_array.tag0\[3\]\[20\] _03748_
+ VGND VGND VPWR VPWR _03749_ sky130_fd_sc_hd__a221o_1
XFILLER_179_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07394_ net1628 _04633_ _04637_ net1202 VGND VGND VPWR VPWR _04640_ sky130_fd_sc_hd__a22o_1
XFILLER_148_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09133_ net1010 net3381 net566 VGND VGND VPWR VPWR _00887_ sky130_fd_sc_hd__mux2_1
X_06345_ tag_array.tag0\[13\]\[14\] net1559 net1463 tag_array.tag0\[14\]\[14\] VGND
+ VGND VPWR VPWR _03686_ sky130_fd_sc_hd__a22o_1
XFILLER_163_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09064_ net1028 net3089 net416 VGND VGND VPWR VPWR _00818_ sky130_fd_sc_hd__mux2_1
X_06276_ tag_array.tag0\[8\]\[8\] net1410 net1316 tag_array.tag0\[11\]\[8\] _03622_
+ VGND VGND VPWR VPWR _03623_ sky130_fd_sc_hd__a221o_1
XFILLER_175_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08015_ data_array.data1\[5\]\[52\] net1545 net1449 data_array.data1\[6\]\[52\] VGND
+ VGND VPWR VPWR _05204_ sky130_fd_sc_hd__a22o_1
XFILLER_163_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold620 data_array.data1\[0\]\[63\] VGND VGND VPWR VPWR net2271 sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 data_array.data0\[1\]\[30\] VGND VGND VPWR VPWR net2282 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold642 tag_array.tag0\[11\]\[2\] VGND VGND VPWR VPWR net2293 sky130_fd_sc_hd__dlygate4sd3_1
Xhold653 data_array.data1\[1\]\[16\] VGND VGND VPWR VPWR net2304 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold664 data_array.data1\[4\]\[53\] VGND VGND VPWR VPWR net2315 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold675 data_array.data0\[4\]\[25\] VGND VGND VPWR VPWR net2326 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold686 data_array.data0\[11\]\[62\] VGND VGND VPWR VPWR net2337 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold697 data_array.data0\[0\]\[33\] VGND VGND VPWR VPWR net2348 sky130_fd_sc_hd__dlygate4sd3_1
X_09966_ net964 net2910 net377 VGND VGND VPWR VPWR _01715_ sky130_fd_sc_hd__mux2_1
Xhold2010 tag_array.tag1\[3\]\[7\] VGND VGND VPWR VPWR net3661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2021 tag_array.tag1\[6\]\[11\] VGND VGND VPWR VPWR net3672 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2032 data_array.data0\[12\]\[57\] VGND VGND VPWR VPWR net3683 sky130_fd_sc_hd__dlygate4sd3_1
X_08917_ net1096 net2942 net431 VGND VGND VPWR VPWR _00673_ sky130_fd_sc_hd__mux2_1
XFILLER_76_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2043 data_array.data0\[9\]\[10\] VGND VGND VPWR VPWR net3694 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2054 data_array.data0\[15\]\[19\] VGND VGND VPWR VPWR net3705 sky130_fd_sc_hd__dlygate4sd3_1
X_09897_ net880 net3742 net381 VGND VGND VPWR VPWR _01647_ sky130_fd_sc_hd__mux2_1
Xhold2065 tag_array.tag1\[9\]\[9\] VGND VGND VPWR VPWR net3716 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1320 data_array.data1\[4\]\[54\] VGND VGND VPWR VPWR net2971 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_96_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_96_clk sky130_fd_sc_hd__clkbuf_8
Xhold1331 data_array.data1\[5\]\[34\] VGND VGND VPWR VPWR net2982 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2076 data_array.data0\[14\]\[36\] VGND VGND VPWR VPWR net3727 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2087 data_array.data1\[7\]\[33\] VGND VGND VPWR VPWR net3738 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1342 tag_array.tag0\[10\]\[18\] VGND VGND VPWR VPWR net2993 sky130_fd_sc_hd__dlygate4sd3_1
X_08848_ _05361_ _05414_ VGND VGND VPWR VPWR _05608_ sky130_fd_sc_hd__or2_1
Xhold1353 data_array.data0\[0\]\[54\] VGND VGND VPWR VPWR net3004 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2098 data_array.data0\[9\]\[34\] VGND VGND VPWR VPWR net3749 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1364 data_array.data1\[13\]\[60\] VGND VGND VPWR VPWR net3015 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1375 data_array.data0\[6\]\[35\] VGND VGND VPWR VPWR net3026 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1386 data_array.data1\[5\]\[35\] VGND VGND VPWR VPWR net3037 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1397 data_array.data1\[12\]\[61\] VGND VGND VPWR VPWR net3048 sky130_fd_sc_hd__dlygate4sd3_1
X_08779_ net709 net2597 net451 VGND VGND VPWR VPWR _00538_ sky130_fd_sc_hd__mux2_1
X_10810_ net2299 net990 net508 VGND VGND VPWR VPWR _02555_ sky130_fd_sc_hd__mux2_1
X_11790_ clknet_leaf_12_clk _00598_ VGND VGND VPWR VPWR data_array.data0\[8\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_0_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_936 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10741_ net1008 net4617 net490 VGND VGND VPWR VPWR _02486_ sky130_fd_sc_hd__mux2_1
X_13460_ clknet_leaf_157_clk _02090_ VGND VGND VPWR VPWR tag_array.tag0\[1\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_10672_ net1875 net1030 net487 VGND VGND VPWR VPWR _02417_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12411_ clknet_leaf_54_clk _01105_ VGND VGND VPWR VPWR data_array.data0\[14\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_97_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13391_ clknet_leaf_34_clk _02021_ VGND VGND VPWR VPWR data_array.data1\[8\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_20_clk clknet_5_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_8
X_12342_ clknet_leaf_80_clk _00016_ VGND VGND VPWR VPWR data_array.rdata0\[24\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_58_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12273_ clknet_leaf_136_clk _01031_ VGND VGND VPWR VPWR tag_array.tag1\[13\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_75_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14012_ clknet_leaf_212_clk _02641_ VGND VGND VPWR VPWR data_array.data1\[5\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
X_11224_ net878 net2998 net652 VGND VGND VPWR VPWR _02967_ sky130_fd_sc_hd__mux2_1
XFILLER_4_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_1023 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11155_ net899 net3717 net541 VGND VGND VPWR VPWR _02898_ sky130_fd_sc_hd__mux2_1
XFILLER_122_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10106_ net2676 net700 net643 VGND VGND VPWR VPWR _01855_ sky130_fd_sc_hd__mux2_1
XFILLER_110_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11086_ net3021 net916 net334 VGND VGND VPWR VPWR _02829_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_87_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_87_clk sky130_fd_sc_hd__clkbuf_8
X_10037_ net938 net2422 net561 VGND VGND VPWR VPWR _01786_ sky130_fd_sc_hd__mux2_1
XFILLER_64_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_19_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11988_ clknet_leaf_109_clk _00796_ VGND VGND VPWR VPWR data_array.data0\[4\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13727_ clknet_leaf_200_clk _02356_ VGND VGND VPWR VPWR data_array.data1\[1\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_10939_ net984 net4389 net531 VGND VGND VPWR VPWR _02684_ sky130_fd_sc_hd__mux2_1
XFILLER_143_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_154_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13658_ clknet_leaf_46_clk _02287_ VGND VGND VPWR VPWR data_array.data1\[15\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_158_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12609_ clknet_leaf_157_clk _01303_ VGND VGND VPWR VPWR tag_array.tag0\[0\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_171_3654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13589_ clknet_leaf_50_clk _02218_ VGND VGND VPWR VPWR data_array.data0\[9\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_11_clk clknet_5_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_30_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06130_ data_array.rdata0\[45\] net1138 net1113 data_array.rdata1\[45\] VGND VGND
+ VPWR VPWR net302 sky130_fd_sc_hd__a22o_1
XFILLER_129_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06061_ net1163 net13 fsm.tag_out1\[13\] net1132 VGND VGND VPWR VPWR _03494_ sky130_fd_sc_hd__a22o_1
XFILLER_133_808 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout407 net408 VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__buf_4
X_09820_ net928 net2521 net387 VGND VGND VPWR VPWR _01571_ sky130_fd_sc_hd__mux2_1
Xfanout418 net425 VGND VGND VPWR VPWR net418 sky130_fd_sc_hd__clkbuf_8
Xfanout429 net433 VGND VGND VPWR VPWR net429 sky130_fd_sc_hd__buf_4
XFILLER_101_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09751_ net1845 net782 net666 VGND VGND VPWR VPWR _01503_ sky130_fd_sc_hd__mux2_1
X_06963_ data_array.data0\[1\]\[20\] net1603 net1507 data_array.data0\[2\]\[20\] VGND
+ VGND VPWR VPWR _04248_ sky130_fd_sc_hd__a22o_1
XFILLER_39_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_78_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_78_clk sky130_fd_sc_hd__clkbuf_8
X_08702_ net2880 net714 net488 VGND VGND VPWR VPWR _00461_ sky130_fd_sc_hd__mux2_1
X_05914_ net118 net1152 _03402_ _03403_ VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__a22o_1
X_09682_ net758 net4524 net607 VGND VGND VPWR VPWR _01434_ sky130_fd_sc_hd__mux2_1
X_06894_ data_array.data0\[4\]\[14\] net1379 net1285 data_array.data0\[7\]\[14\] _04184_
+ VGND VGND VPWR VPWR _04185_ sky130_fd_sc_hd__a221o_1
X_08633_ net1923 net791 net507 VGND VGND VPWR VPWR _00392_ sky130_fd_sc_hd__mux2_1
X_05845_ net143 net1155 _03356_ _03357_ VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__a22o_1
XFILLER_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08564_ net700 net4300 net589 VGND VGND VPWR VPWR _00332_ sky130_fd_sc_hd__mux2_1
XFILLER_54_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05776_ _03291_ _03292_ _03263_ _03266_ VGND VGND VPWR VPWR _03293_ sky130_fd_sc_hd__a211o_1
XFILLER_70_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07515_ net1614 _04743_ _04747_ net1188 VGND VGND VPWR VPWR _04750_ sky130_fd_sc_hd__a22o_1
X_08495_ net822 net813 net854 _05547_ VGND VGND VPWR VPWR _05567_ sky130_fd_sc_hd__or4b_4
X_07446_ data_array.data1\[8\]\[0\] net1366 net1272 data_array.data1\[11\]\[0\] _04686_
+ VGND VGND VPWR VPWR _04687_ sky130_fd_sc_hd__a221o_1
XFILLER_22_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_963 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07377_ data_array.data0\[5\]\[58\] net1546 net1450 data_array.data0\[6\]\[58\] VGND
+ VGND VPWR VPWR _04624_ sky130_fd_sc_hd__a22o_1
XFILLER_10_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09116_ net1079 net3941 net568 VGND VGND VPWR VPWR _00870_ sky130_fd_sc_hd__mux2_1
XFILLER_164_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06328_ net1182 _03665_ _03669_ net1230 VGND VGND VPWR VPWR _03671_ sky130_fd_sc_hd__a22o_1
XFILLER_163_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09047_ net1096 net4228 net415 VGND VGND VPWR VPWR _00801_ sky130_fd_sc_hd__mux2_1
X_06259_ tag_array.tag0\[1\]\[6\] net1564 net1468 tag_array.tag0\[2\]\[6\] VGND VGND
+ VPWR VPWR _03608_ sky130_fd_sc_hd__a22o_1
XFILLER_163_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_92_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold450 data_array.data1\[0\]\[60\] VGND VGND VPWR VPWR net2101 sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 data_array.data1\[10\]\[13\] VGND VGND VPWR VPWR net2112 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold472 tag_array.tag1\[14\]\[24\] VGND VGND VPWR VPWR net2123 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold483 data_array.data0\[4\]\[12\] VGND VGND VPWR VPWR net2134 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold494 data_array.data1\[1\]\[31\] VGND VGND VPWR VPWR net2145 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_70_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout930 _05510_ VGND VGND VPWR VPWR net930 sky130_fd_sc_hd__clkbuf_2
Xfanout941 _05504_ VGND VGND VPWR VPWR net941 sky130_fd_sc_hd__dlymetal6s2s_1
X_09949_ net1033 net3222 net375 VGND VGND VPWR VPWR _01698_ sky130_fd_sc_hd__mux2_1
Xfanout952 _05498_ VGND VGND VPWR VPWR net952 sky130_fd_sc_hd__clkbuf_2
XFILLER_49_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout963 _05494_ VGND VGND VPWR VPWR net963 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_69_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_69_clk sky130_fd_sc_hd__clkbuf_8
Xfanout974 _05488_ VGND VGND VPWR VPWR net974 sky130_fd_sc_hd__clkbuf_2
Xfanout985 _05482_ VGND VGND VPWR VPWR net985 sky130_fd_sc_hd__buf_1
Xfanout996 net999 VGND VGND VPWR VPWR net996 sky130_fd_sc_hd__clkbuf_2
X_12960_ clknet_leaf_106_clk _01654_ VGND VGND VPWR VPWR tag_array.tag0\[4\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_180_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1150 data_array.data0\[5\]\[45\] VGND VGND VPWR VPWR net2801 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1161 tag_array.tag0\[4\]\[17\] VGND VGND VPWR VPWR net2812 sky130_fd_sc_hd__dlygate4sd3_1
X_11911_ clknet_leaf_62_clk _00719_ VGND VGND VPWR VPWR data_array.data0\[5\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1172 data_array.data1\[15\]\[19\] VGND VGND VPWR VPWR net2823 sky130_fd_sc_hd__dlygate4sd3_1
X_12891_ clknet_leaf_54_clk _01585_ VGND VGND VPWR VPWR data_array.data0\[12\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1183 tag_array.tag0\[5\]\[23\] VGND VGND VPWR VPWR net2834 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1194 data_array.data1\[6\]\[56\] VGND VGND VPWR VPWR net2845 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11842_ clknet_leaf_87_clk _00650_ VGND VGND VPWR VPWR data_array.data0\[7\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_16_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11773_ clknet_leaf_235_clk _00581_ VGND VGND VPWR VPWR data_array.data0\[8\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13512_ clknet_leaf_58_clk _02141_ VGND VGND VPWR VPWR data_array.data1\[0\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_10724_ net1078 net2673 net492 VGND VGND VPWR VPWR _02469_ sky130_fd_sc_hd__mux2_1
X_14492_ clknet_leaf_161_clk _03115_ VGND VGND VPWR VPWR tag_array.dirty0\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_158_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13443_ clknet_leaf_193_clk _02073_ VGND VGND VPWR VPWR data_array.data1\[8\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10655_ net2060 net1098 net483 VGND VGND VPWR VPWR _02400_ sky130_fd_sc_hd__mux2_1
XFILLER_16_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload17 clknet_leaf_2_clk VGND VGND VPWR VPWR clkload17/Y sky130_fd_sc_hd__clkinv_4
XFILLER_103_1044 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13374_ clknet_leaf_102_clk _02004_ VGND VGND VPWR VPWR tag_array.tag0\[2\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_10586_ net862 net3121 net463 VGND VGND VPWR VPWR _02331_ sky130_fd_sc_hd__mux2_1
Xclkload28 clknet_leaf_267_clk VGND VGND VPWR VPWR clkload28/Y sky130_fd_sc_hd__inv_6
Xclkload39 clknet_leaf_18_clk VGND VGND VPWR VPWR clkload39/Y sky130_fd_sc_hd__bufinv_16
X_12325_ clknet_leaf_81_clk _00061_ VGND VGND VPWR VPWR data_array.rdata0\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_103_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_454 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12256_ clknet_leaf_134_clk _01014_ VGND VGND VPWR VPWR tag_array.tag1\[14\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_108_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11207_ net947 net4421 net648 VGND VGND VPWR VPWR _02950_ sky130_fd_sc_hd__mux2_1
X_12187_ clknet_leaf_160_clk _00995_ VGND VGND VPWR VPWR tag_array.tag0\[14\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_68_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11138_ net966 net3850 net549 VGND VGND VPWR VPWR _02881_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_147_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_6__f_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_5_6__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_68_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_147_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11069_ net2514 net986 net334 VGND VGND VPWR VPWR _02812_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_0_clk clknet_5_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_37_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05630_ fsm.lru_out dirty_way0 fsm.valid0 VGND VGND VPWR VPWR _03149_ sky130_fd_sc_hd__and3b_1
XFILLER_92_997 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07300_ data_array.data0\[5\]\[51\] net1522 net1426 data_array.data0\[6\]\[51\] VGND
+ VGND VPWR VPWR _04554_ sky130_fd_sc_hd__a22o_1
X_08280_ net121 net56 net1639 VGND VGND VPWR VPWR _05423_ sky130_fd_sc_hd__mux2_1
XFILLER_20_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07231_ _04490_ _04491_ VGND VGND VPWR VPWR _00038_ sky130_fd_sc_hd__or2_1
XFILLER_118_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07162_ data_array.data0\[4\]\[38\] net1396 net1302 data_array.data0\[7\]\[38\] _04428_
+ VGND VGND VPWR VPWR _04429_ sky130_fd_sc_hd__a221o_1
XFILLER_145_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06113_ data_array.rdata0\[28\] net1135 net1112 data_array.rdata1\[28\] VGND VGND
+ VPWR VPWR net283 sky130_fd_sc_hd__a22o_1
X_07093_ data_array.data0\[9\]\[32\] net1523 net1427 data_array.data0\[10\]\[32\]
+ VGND VGND VPWR VPWR _04366_ sky130_fd_sc_hd__a22o_1
XFILLER_172_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06044_ fsm.tag_out0\[4\] net1120 _03485_ VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__a21o_1
XFILLER_132_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09803_ net998 net4603 net390 VGND VGND VPWR VPWR _01554_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_184_3889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07995_ data_array.data1\[13\]\[50\] net1527 net1431 data_array.data1\[14\]\[50\]
+ VGND VGND VPWR VPWR _05186_ sky130_fd_sc_hd__a22o_1
X_09734_ net751 net2456 net684 VGND VGND VPWR VPWR _01486_ sky130_fd_sc_hd__mux2_1
X_06946_ data_array.data0\[13\]\[19\] net1582 net1486 data_array.data0\[14\]\[19\]
+ VGND VGND VPWR VPWR _04232_ sky130_fd_sc_hd__a22o_1
XFILLER_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09665_ net727 net4598 net613 VGND VGND VPWR VPWR _01417_ sky130_fd_sc_hd__mux2_1
X_06877_ net1629 _04163_ _04167_ net1203 VGND VGND VPWR VPWR _04170_ sky130_fd_sc_hd__a22o_1
XFILLER_28_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08616_ net759 net2915 net524 VGND VGND VPWR VPWR _00375_ sky130_fd_sc_hd__mux2_1
XFILLER_82_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05828_ _03274_ _03283_ fsm.valid1 VGND VGND VPWR VPWR _03345_ sky130_fd_sc_hd__or3b_1
X_09596_ net965 net4262 net400 VGND VGND VPWR VPWR _01348_ sky130_fd_sc_hd__mux2_1
XFILLER_42_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08547_ net766 net4581 net583 VGND VGND VPWR VPWR _00315_ sky130_fd_sc_hd__mux2_1
X_05759_ net20 _03144_ _03269_ _03270_ _03275_ VGND VGND VPWR VPWR _03276_ sky130_fd_sc_hd__a2111o_1
XFILLER_126_1000 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08478_ net1704 net647 VGND VGND VPWR VPWR _00288_ sky130_fd_sc_hd__nand2b_1
X_07429_ _04670_ _04671_ VGND VGND VPWR VPWR _00058_ sky130_fd_sc_hd__or2_1
XFILLER_24_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_516 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10440_ net3033 net892 net664 VGND VGND VPWR VPWR _02186_ sky130_fd_sc_hd__mux2_1
XFILLER_136_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10371_ net716 net3389 net539 VGND VGND VPWR VPWR _02118_ sky130_fd_sc_hd__mux2_1
XFILLER_152_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12110_ clknet_leaf_21_clk _00918_ VGND VGND VPWR VPWR data_array.data1\[14\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13090_ clknet_leaf_258_clk _01784_ VGND VGND VPWR VPWR data_array.data1\[13\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_152_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12041_ clknet_leaf_1_clk _00849_ VGND VGND VPWR VPWR data_array.data0\[6\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_979 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold280 data_array.data0\[0\]\[1\] VGND VGND VPWR VPWR net1931 sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 data_array.data1\[1\]\[36\] VGND VGND VPWR VPWR net1942 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout760 net761 VGND VGND VPWR VPWR net760 sky130_fd_sc_hd__clkbuf_2
Xfanout771 _05375_ VGND VGND VPWR VPWR net771 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout782 _05369_ VGND VGND VPWR VPWR net782 sky130_fd_sc_hd__clkbuf_2
XFILLER_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13992_ clknet_leaf_265_clk _02621_ VGND VGND VPWR VPWR data_array.data1\[5\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout793 _05365_ VGND VGND VPWR VPWR net793 sky130_fd_sc_hd__clkbuf_2
X_12943_ clknet_leaf_38_clk _01637_ VGND VGND VPWR VPWR data_array.data0\[13\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_65_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_142_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12874_ clknet_leaf_87_clk _01568_ VGND VGND VPWR VPWR data_array.data0\[12\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_46_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11825_ clknet_leaf_229_clk _00633_ VGND VGND VPWR VPWR data_array.data0\[7\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_103_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11756_ clknet_leaf_22_clk _00564_ VGND VGND VPWR VPWR data_array.data0\[8\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_120_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10707_ net3992 net890 net479 VGND VGND VPWR VPWR _02452_ sky130_fd_sc_hd__mux2_1
X_14475_ clknet_leaf_55_clk _03098_ VGND VGND VPWR VPWR data_array.data1\[7\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
X_11687_ clknet_leaf_191_clk _00495_ VGND VGND VPWR VPWR tag_array.tag1\[15\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_13426_ clknet_leaf_244_clk _02056_ VGND VGND VPWR VPWR data_array.data1\[8\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
X_10638_ net1847 net908 net466 VGND VGND VPWR VPWR _02383_ sky130_fd_sc_hd__mux2_1
Xclkload106 clknet_leaf_91_clk VGND VGND VPWR VPWR clkload106/X sky130_fd_sc_hd__clkbuf_8
Xclkload117 clknet_leaf_73_clk VGND VGND VPWR VPWR clkload117/X sky130_fd_sc_hd__clkbuf_8
Xclkload128 clknet_leaf_83_clk VGND VGND VPWR VPWR clkload128/Y sky130_fd_sc_hd__inv_6
Xclkload139 clknet_leaf_221_clk VGND VGND VPWR VPWR clkload139/X sky130_fd_sc_hd__clkbuf_8
XFILLER_60_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13357_ clknet_leaf_168_clk _01987_ VGND VGND VPWR VPWR tag_array.tag0\[2\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_10569_ net930 net3054 net455 VGND VGND VPWR VPWR _02314_ sky130_fd_sc_hd__mux2_1
X_12308_ clknet_leaf_100_clk _01066_ VGND VGND VPWR VPWR tag_array.tag1\[12\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_154_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13288_ clknet_leaf_192_clk _01918_ VGND VGND VPWR VPWR data_array.data0\[11\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
X_12239_ clknet_leaf_151_clk _00169_ VGND VGND VPWR VPWR fsm.tag_out1\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_170_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_166_3553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2609 data_array.data0\[7\]\[40\] VGND VGND VPWR VPWR net4260 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_127_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1908 data_array.data1\[11\]\[63\] VGND VGND VPWR VPWR net3559 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_110_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06800_ net1622 _04093_ _04097_ net1196 VGND VGND VPWR VPWR _04100_ sky130_fd_sc_hd__a22o_1
Xhold1919 data_array.data1\[15\]\[2\] VGND VGND VPWR VPWR net3570 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_110_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07780_ net1178 _04985_ _04989_ net1226 VGND VGND VPWR VPWR _04991_ sky130_fd_sc_hd__a22o_1
XFILLER_7_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput4 cpu_addr[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_2
XFILLER_65_931 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06731_ tag_array.tag1\[8\]\[24\] net1372 net1278 tag_array.tag1\[11\]\[24\] _04036_
+ VGND VGND VPWR VPWR _04037_ sky130_fd_sc_hd__a221o_1
XFILLER_36_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09450_ net864 net3499 net582 VGND VGND VPWR VPWR _01203_ sky130_fd_sc_hd__mux2_1
XFILLER_149_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06662_ tag_array.tag1\[1\]\[18\] net1562 net1466 tag_array.tag1\[2\]\[18\] VGND
+ VGND VPWR VPWR _03974_ sky130_fd_sc_hd__a22o_1
XFILLER_24_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08401_ net1130 _05503_ VGND VGND VPWR VPWR _05504_ sky130_fd_sc_hd__and2_1
XFILLER_36_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05613_ net31 VGND VGND VPWR VPWR _03135_ sky130_fd_sc_hd__inv_2
X_09381_ net877 net3855 net405 VGND VGND VPWR VPWR _01134_ sky130_fd_sc_hd__mux2_1
X_06593_ _03910_ _03911_ VGND VGND VPWR VPWR _00158_ sky130_fd_sc_hd__or2_2
X_08332_ net1127 _05457_ VGND VGND VPWR VPWR _05458_ sky130_fd_sc_hd__and2_1
XFILLER_32_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08263_ net1650 net1164 net24 VGND VGND VPWR VPWR _05410_ sky130_fd_sc_hd__and3_1
X_07214_ data_array.data0\[13\]\[43\] net1569 net1473 data_array.data0\[14\]\[43\]
+ VGND VGND VPWR VPWR _04476_ sky130_fd_sc_hd__a22o_1
X_08194_ fsm.state\[2\] net1644 net840 VGND VGND VPWR VPWR _05364_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_41_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07145_ data_array.data0\[8\]\[37\] net1356 net1262 data_array.data0\[11\]\[37\]
+ _04412_ VGND VGND VPWR VPWR _04413_ sky130_fd_sc_hd__a221o_1
XFILLER_119_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07076_ net1178 _04345_ _04349_ net1226 VGND VGND VPWR VPWR _04351_ sky130_fd_sc_hd__a22o_1
XFILLER_156_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06027_ fsm.lru_out fsm.state\[5\] fsm.valid0 VGND VGND VPWR VPWR _03477_ sky130_fd_sc_hd__and3b_4
XTAP_TAPCELL_ROW_7_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_184_Left_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07978_ net1179 _05165_ _05169_ net1227 VGND VGND VPWR VPWR _05171_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_87_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09717_ net720 net2684 net609 VGND VGND VPWR VPWR _01469_ sky130_fd_sc_hd__mux2_1
X_06929_ data_array.data0\[8\]\[17\] net1339 net1245 data_array.data0\[11\]\[17\]
+ _04216_ VGND VGND VPWR VPWR _04217_ sky130_fd_sc_hd__a221o_1
XFILLER_132_1070 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09648_ net697 net3637 net615 VGND VGND VPWR VPWR _01400_ sky130_fd_sc_hd__mux2_1
XFILLER_27_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09579_ net1033 net3705 net399 VGND VGND VPWR VPWR _01331_ sky130_fd_sc_hd__mux2_1
XFILLER_35_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11610_ clknet_leaf_99_clk _00418_ VGND VGND VPWR VPWR tag_array.tag1\[3\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_26_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12590_ clknet_leaf_186_clk _01284_ VGND VGND VPWR VPWR tag_array.tag0\[10\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_143_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11541_ clknet_leaf_129_clk _00349_ VGND VGND VPWR VPWR tag_array.tag1\[6\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14260_ clknet_leaf_79_clk _02889_ VGND VGND VPWR VPWR data_array.data1\[12\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11472_ clknet_leaf_206_clk _00282_ VGND VGND VPWR VPWR data_array.data0\[0\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13211_ clknet_leaf_76_clk _00106_ VGND VGND VPWR VPWR data_array.rdata1\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10423_ net3577 net963 net664 VGND VGND VPWR VPWR _02169_ sky130_fd_sc_hd__mux2_1
X_14191_ clknet_leaf_235_clk _02820_ VGND VGND VPWR VPWR data_array.data0\[2\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_100_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13142_ clknet_leaf_196_clk _01836_ VGND VGND VPWR VPWR tag_array.tag1\[8\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_10354_ net785 net2760 net538 VGND VGND VPWR VPWR _02101_ sky130_fd_sc_hd__mux2_1
XFILLER_83_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13073_ clknet_leaf_93_clk _01767_ VGND VGND VPWR VPWR data_array.data1\[13\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10285_ net2195 net1021 net635 VGND VGND VPWR VPWR _02032_ sky130_fd_sc_hd__mux2_1
X_12024_ clknet_leaf_11_clk _00832_ VGND VGND VPWR VPWR data_array.data0\[6\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout1500 net1517 VGND VGND VPWR VPWR net1500 sky130_fd_sc_hd__clkbuf_4
Xfanout1511 net1513 VGND VGND VPWR VPWR net1511 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_168_Right_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1522 net1524 VGND VGND VPWR VPWR net1522 sky130_fd_sc_hd__clkbuf_4
XFILLER_78_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1533 net1543 VGND VGND VPWR VPWR net1533 sky130_fd_sc_hd__buf_2
XFILLER_78_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_144_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1544 net1546 VGND VGND VPWR VPWR net1544 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_144_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1555 net1557 VGND VGND VPWR VPWR net1555 sky130_fd_sc_hd__clkbuf_4
XFILLER_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1566 _03508_ VGND VGND VPWR VPWR net1566 sky130_fd_sc_hd__buf_2
Xfanout1577 net1579 VGND VGND VPWR VPWR net1577 sky130_fd_sc_hd__clkbuf_4
Xfanout1588 net1590 VGND VGND VPWR VPWR net1588 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_161_3450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout590 _05591_ VGND VGND VPWR VPWR net590 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_161_3461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1599 net1600 VGND VGND VPWR VPWR net1599 sky130_fd_sc_hd__buf_2
X_13975_ clknet_leaf_64_clk _02604_ VGND VGND VPWR VPWR data_array.data1\[5\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_46_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12926_ clknet_leaf_71_clk _01620_ VGND VGND VPWR VPWR data_array.data0\[13\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12857_ clknet_leaf_262_clk _01551_ VGND VGND VPWR VPWR data_array.data0\[12\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11808_ clknet_leaf_111_clk _00616_ VGND VGND VPWR VPWR data_array.data0\[7\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_12788_ clknet_leaf_195_clk _01482_ VGND VGND VPWR VPWR tag_array.tag1\[10\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_11739_ clknet_leaf_204_clk _00547_ VGND VGND VPWR VPWR data_array.data0\[8\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_14458_ clknet_leaf_87_clk _03081_ VGND VGND VPWR VPWR data_array.data1\[7\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_174_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13409_ clknet_leaf_39_clk _02039_ VGND VGND VPWR VPWR data_array.data1\[8\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_14389_ clknet_leaf_240_clk _03012_ VGND VGND VPWR VPWR data_array.data1\[10\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_170_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08950_ net964 net2498 net432 VGND VGND VPWR VPWR _00706_ sky130_fd_sc_hd__mux2_1
X_07901_ net1166 _05095_ _05099_ net1214 VGND VGND VPWR VPWR _05101_ sky130_fd_sc_hd__a22o_1
Xhold2406 data_array.data0\[3\]\[34\] VGND VGND VPWR VPWR net4057 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08881_ net982 net4195 net434 VGND VGND VPWR VPWR _00638_ sky130_fd_sc_hd__mux2_1
Xhold2417 data_array.data0\[10\]\[18\] VGND VGND VPWR VPWR net4068 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_181_3837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2428 data_array.data1\[3\]\[11\] VGND VGND VPWR VPWR net4079 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_135_Right_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2439 lru_array.lru_mem\[0\] VGND VGND VPWR VPWR net4090 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_5_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1705 data_array.data1\[12\]\[21\] VGND VGND VPWR VPWR net3356 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1716 data_array.data0\[12\]\[30\] VGND VGND VPWR VPWR net3367 sky130_fd_sc_hd__dlygate4sd3_1
X_07832_ data_array.data1\[1\]\[35\] net1525 net1429 data_array.data1\[2\]\[35\] VGND
+ VGND VPWR VPWR _05038_ sky130_fd_sc_hd__a22o_1
XFILLER_29_419 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1727 tag_array.tag1\[13\]\[19\] VGND VGND VPWR VPWR net3378 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1738 tag_array.tag0\[15\]\[19\] VGND VGND VPWR VPWR net3389 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1749 data_array.data0\[3\]\[43\] VGND VGND VPWR VPWR net3400 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_110_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07763_ data_array.data1\[0\]\[29\] net1381 net1287 data_array.data1\[3\]\[29\] _04974_
+ VGND VGND VPWR VPWR _04975_ sky130_fd_sc_hd__a221o_1
X_09502_ net719 net3155 net624 VGND VGND VPWR VPWR _01255_ sky130_fd_sc_hd__mux2_1
X_06714_ _04020_ _04021_ VGND VGND VPWR VPWR _00170_ sky130_fd_sc_hd__or2_1
XFILLER_71_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07694_ data_array.data1\[13\]\[23\] net1550 net1454 data_array.data1\[14\]\[23\]
+ VGND VGND VPWR VPWR _04912_ sky130_fd_sc_hd__a22o_1
XFILLER_80_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09433_ net934 net3295 net587 VGND VGND VPWR VPWR _01186_ sky130_fd_sc_hd__mux2_1
X_06645_ tag_array.tag1\[4\]\[16\] net1417 net1323 tag_array.tag1\[7\]\[16\] _03958_
+ VGND VGND VPWR VPWR _03959_ sky130_fd_sc_hd__a221o_1
XFILLER_24_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_179_3799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09364_ net945 net3062 net402 VGND VGND VPWR VPWR _01117_ sky130_fd_sc_hd__mux2_1
XFILLER_80_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06576_ tag_array.tag1\[9\]\[10\] net1595 net1499 tag_array.tag1\[10\]\[10\] VGND
+ VGND VPWR VPWR _03896_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_23_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08315_ net2384 net1058 net688 VGND VGND VPWR VPWR _00234_ sky130_fd_sc_hd__mux2_1
XFILLER_178_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09295_ net701 net3745 net564 VGND VGND VPWR VPWR _01049_ sky130_fd_sc_hd__mux2_1
XANTENNA_20 _03506_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_31 net331 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_42 net518 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_53 net1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08246_ fsm.tag_out1\[17\] net817 net809 fsm.tag_out0\[17\] _05398_ VGND VGND VPWR
+ VPWR _05399_ sky130_fd_sc_hd__a221o_2
XFILLER_21_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_64 net1613 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_75 _05385_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_86 net1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08177_ _05350_ _05351_ VGND VGND VPWR VPWR _00128_ sky130_fd_sc_hd__or2_1
XFILLER_118_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07128_ data_array.data0\[1\]\[35\] net1527 net1431 data_array.data0\[2\]\[35\] VGND
+ VGND VPWR VPWR _04398_ sky130_fd_sc_hd__a22o_1
XFILLER_107_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07059_ data_array.data0\[0\]\[29\] net1379 net1285 data_array.data0\[3\]\[29\] _04334_
+ VGND VGND VPWR VPWR _04335_ sky130_fd_sc_hd__a221o_1
Xoutput171 net171 VGND VGND VPWR VPWR cpu_rdata[15] sky130_fd_sc_hd__buf_6
Xoutput182 net182 VGND VGND VPWR VPWR cpu_rdata[25] sky130_fd_sc_hd__buf_4
XFILLER_153_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput193 net193 VGND VGND VPWR VPWR cpu_rdata[35] sky130_fd_sc_hd__buf_4
X_10070_ net745 net3737 net599 VGND VGND VPWR VPWR _01819_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_102_Right_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2940 data_array.data0\[7\]\[57\] VGND VGND VPWR VPWR net4591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2951 data_array.data0\[14\]\[1\] VGND VGND VPWR VPWR net4602 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2962 tag_array.tag1\[6\]\[20\] VGND VGND VPWR VPWR net4613 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2973 fsm.state\[0\] VGND VGND VPWR VPWR net4624 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_986 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13760_ clknet_leaf_9_clk _02389_ VGND VGND VPWR VPWR data_array.data1\[1\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_44_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10972_ net807 _05587_ VGND VGND VPWR VPWR _03132_ sky130_fd_sc_hd__and2_4
XFILLER_83_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12711_ clknet_leaf_178_clk _01405_ VGND VGND VPWR VPWR tag_array.tag0\[7\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_13691_ clknet_leaf_4_clk _02320_ VGND VGND VPWR VPWR data_array.data1\[15\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_44_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12642_ clknet_leaf_97_clk _01336_ VGND VGND VPWR VPWR data_array.data0\[15\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12573_ clknet_leaf_138_clk _01267_ VGND VGND VPWR VPWR tag_array.tag0\[10\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_178_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11524_ clknet_leaf_130_clk _00332_ VGND VGND VPWR VPWR tag_array.tag1\[9\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_14312_ clknet_leaf_257_clk _02941_ VGND VGND VPWR VPWR data_array.data1\[11\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14243_ clknet_leaf_221_clk _02872_ VGND VGND VPWR VPWR data_array.data1\[12\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11455_ clknet_leaf_86_clk _00265_ VGND VGND VPWR VPWR data_array.data0\[0\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_125_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10406_ net2820 net1030 net671 VGND VGND VPWR VPWR _02152_ sky130_fd_sc_hd__mux2_1
Xclkbuf_5_31__f_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_5_31__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_14174_ clknet_leaf_8_clk _02803_ VGND VGND VPWR VPWR data_array.data0\[2\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_78_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11386_ clknet_leaf_97_clk _00196_ VGND VGND VPWR VPWR tag_array.tag1\[7\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_152_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13125_ clknet_leaf_163_clk _01819_ VGND VGND VPWR VPWR tag_array.tag0\[3\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_10337_ net751 net3864 net592 VGND VGND VPWR VPWR _02084_ sky130_fd_sc_hd__mux2_1
XFILLER_139_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_163_3501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ clknet_leaf_82_clk _01750_ VGND VGND VPWR VPWR data_array.data1\[13\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10268_ net2031 net1090 net637 VGND VGND VPWR VPWR _02015_ sky130_fd_sc_hd__mux2_1
X_12007_ clknet_leaf_249_clk _00815_ VGND VGND VPWR VPWR data_array.data0\[6\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout1330 net1331 VGND VGND VPWR VPWR net1330 sky130_fd_sc_hd__clkbuf_4
Xfanout1341 net1342 VGND VGND VPWR VPWR net1341 sky130_fd_sc_hd__clkbuf_4
Xfanout1352 net1376 VGND VGND VPWR VPWR net1352 sky130_fd_sc_hd__buf_2
X_10199_ net1009 net3718 net354 VGND VGND VPWR VPWR _01946_ sky130_fd_sc_hd__mux2_1
Xfanout1363 net1364 VGND VGND VPWR VPWR net1363 sky130_fd_sc_hd__clkbuf_2
Xfanout1374 net1375 VGND VGND VPWR VPWR net1374 sky130_fd_sc_hd__buf_2
Xfanout1385 net1388 VGND VGND VPWR VPWR net1385 sky130_fd_sc_hd__clkbuf_4
XFILLER_94_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1396 net1399 VGND VGND VPWR VPWR net1396 sky130_fd_sc_hd__clkbuf_4
XFILLER_93_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13958_ clknet_leaf_123_clk _02587_ VGND VGND VPWR VPWR data_array.data1\[4\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_98_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12909_ clknet_leaf_206_clk _01603_ VGND VGND VPWR VPWR data_array.data0\[13\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_13889_ clknet_leaf_248_clk _02518_ VGND VGND VPWR VPWR data_array.data1\[3\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
X_06430_ tag_array.tag0\[8\]\[22\] net1374 net1280 tag_array.tag0\[11\]\[22\] _03762_
+ VGND VGND VPWR VPWR _03763_ sky130_fd_sc_hd__a221o_1
XFILLER_179_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06361_ net1229 _03695_ _03699_ net1181 VGND VGND VPWR VPWR _03701_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_174_3696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08100_ _05280_ _05281_ VGND VGND VPWR VPWR _00118_ sky130_fd_sc_hd__or2_1
XFILLER_148_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09080_ net964 net1958 net416 VGND VGND VPWR VPWR _00834_ sky130_fd_sc_hd__mux2_1
XFILLER_174_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06292_ tag_array.tag0\[5\]\[9\] net1598 net1502 tag_array.tag0\[6\]\[9\] VGND VGND
+ VPWR VPWR _03638_ sky130_fd_sc_hd__a22o_1
X_08031_ data_array.data1\[4\]\[53\] net1332 net1238 data_array.data1\[7\]\[53\] _05218_
+ VGND VGND VPWR VPWR _05219_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_135_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput40 cpu_wdata[15] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_135_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput51 cpu_wdata[25] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_1
Xhold802 data_array.data1\[11\]\[60\] VGND VGND VPWR VPWR net2453 sky130_fd_sc_hd__dlygate4sd3_1
Xinput62 cpu_wdata[35] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_1
Xinput73 cpu_wdata[45] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_1
Xhold813 data_array.data0\[2\]\[16\] VGND VGND VPWR VPWR net2464 sky130_fd_sc_hd__dlygate4sd3_1
Xinput84 cpu_wdata[55] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_1
Xinput95 cpu_wdata[7] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_1
Xhold824 data_array.data0\[8\]\[53\] VGND VGND VPWR VPWR net2475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold835 tag_array.tag1\[4\]\[11\] VGND VGND VPWR VPWR net2486 sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 tag_array.tag1\[12\]\[22\] VGND VGND VPWR VPWR net2497 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold857 data_array.data0\[12\]\[6\] VGND VGND VPWR VPWR net2508 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_264_clk clknet_5_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_264_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_66_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09982_ net902 net3337 net372 VGND VGND VPWR VPWR _01731_ sky130_fd_sc_hd__mux2_1
XFILLER_107_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold868 data_array.data0\[7\]\[48\] VGND VGND VPWR VPWR net2519 sky130_fd_sc_hd__dlygate4sd3_1
Xhold879 data_array.data1\[13\]\[52\] VGND VGND VPWR VPWR net2530 sky130_fd_sc_hd__dlygate4sd3_1
X_08933_ net1032 net2473 net430 VGND VGND VPWR VPWR _00689_ sky130_fd_sc_hd__mux2_1
Xhold2203 data_array.data0\[10\]\[4\] VGND VGND VPWR VPWR net3854 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2214 data_array.data0\[13\]\[6\] VGND VGND VPWR VPWR net3865 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2225 data_array.data1\[15\]\[5\] VGND VGND VPWR VPWR net3876 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_36_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2236 data_array.data1\[15\]\[24\] VGND VGND VPWR VPWR net3887 sky130_fd_sc_hd__dlygate4sd3_1
X_08864_ net1048 net3238 net438 VGND VGND VPWR VPWR _00621_ sky130_fd_sc_hd__mux2_1
Xhold2247 data_array.data1\[15\]\[41\] VGND VGND VPWR VPWR net3898 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1502 data_array.data1\[14\]\[11\] VGND VGND VPWR VPWR net3153 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1513 tag_array.tag0\[7\]\[11\] VGND VGND VPWR VPWR net3164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2258 data_array.data0\[7\]\[43\] VGND VGND VPWR VPWR net3909 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1524 data_array.data0\[11\]\[34\] VGND VGND VPWR VPWR net3175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2269 data_array.data1\[3\]\[59\] VGND VGND VPWR VPWR net3920 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1535 tag_array.tag0\[12\]\[15\] VGND VGND VPWR VPWR net3186 sky130_fd_sc_hd__dlygate4sd3_1
X_07815_ data_array.data1\[13\]\[34\] net1532 net1436 data_array.data1\[14\]\[34\]
+ VGND VGND VPWR VPWR _05022_ sky130_fd_sc_hd__a22o_1
XFILLER_96_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1546 data_array.data0\[9\]\[20\] VGND VGND VPWR VPWR net3197 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1557 data_array.data0\[9\]\[18\] VGND VGND VPWR VPWR net3208 sky130_fd_sc_hd__dlygate4sd3_1
X_08795_ net1952 net1065 net446 VGND VGND VPWR VPWR _00553_ sky130_fd_sc_hd__mux2_1
Xhold1568 data_array.data0\[9\]\[41\] VGND VGND VPWR VPWR net3219 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1579 data_array.data0\[5\]\[51\] VGND VGND VPWR VPWR net3230 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_28_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07746_ net1616 _04953_ _04957_ net1191 VGND VGND VPWR VPWR _04960_ sky130_fd_sc_hd__a22o_1
XFILLER_25_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07677_ data_array.data1\[12\]\[21\] net1365 net1271 data_array.data1\[15\]\[21\]
+ _04896_ VGND VGND VPWR VPWR _04897_ sky130_fd_sc_hd__a221o_1
XFILLER_26_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09416_ net1001 net2494 net579 VGND VGND VPWR VPWR _01169_ sky130_fd_sc_hd__mux2_1
XFILLER_52_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06628_ tag_array.tag1\[8\]\[15\] net1401 net1307 tag_array.tag1\[11\]\[15\] _03942_
+ VGND VGND VPWR VPWR _03943_ sky130_fd_sc_hd__a221o_1
X_09347_ net1012 net4532 net406 VGND VGND VPWR VPWR _01100_ sky130_fd_sc_hd__mux2_1
X_06559_ net1184 _03875_ _03879_ net1232 VGND VGND VPWR VPWR _03881_ sky130_fd_sc_hd__a22o_1
XFILLER_32_34 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09278_ net767 net3949 net559 VGND VGND VPWR VPWR _01032_ sky130_fd_sc_hd__mux2_1
XFILLER_138_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08229_ net746 net4210 net800 VGND VGND VPWR VPWR _00207_ sky130_fd_sc_hd__mux2_1
XFILLER_166_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11240_ net1070 net3078 net683 VGND VGND VPWR VPWR _02983_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_95_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_255_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_255_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11171_ net1091 net2506 net652 VGND VGND VPWR VPWR _02914_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10122_ net1059 net3066 net364 VGND VGND VPWR VPWR _01870_ sky130_fd_sc_hd__mux2_1
XFILLER_164_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_983 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10053_ net874 net4013 net561 VGND VGND VPWR VPWR _01802_ sky130_fd_sc_hd__mux2_1
XFILLER_0_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2770 data_array.data1\[11\]\[41\] VGND VGND VPWR VPWR net4421 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2781 data_array.data0\[12\]\[11\] VGND VGND VPWR VPWR net4432 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_36_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2792 data_array.data0\[14\]\[59\] VGND VGND VPWR VPWR net4443 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_180_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13812_ clknet_leaf_83_clk _02441_ VGND VGND VPWR VPWR data_array.data1\[2\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_91_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10955_ _05514_ net3843 net533 VGND VGND VPWR VPWR _02700_ sky130_fd_sc_hd__mux2_1
X_13743_ clknet_leaf_240_clk _02372_ VGND VGND VPWR VPWR data_array.data1\[1\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_139_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13674_ clknet_leaf_7_clk _02303_ VGND VGND VPWR VPWR data_array.data1\[15\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_139_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10886_ net942 net3252 net521 VGND VGND VPWR VPWR _02631_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_156_3360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12625_ clknet_leaf_113_clk _01319_ VGND VGND VPWR VPWR data_array.data0\[15\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_14_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12556_ clknet_leaf_147_clk _01250_ VGND VGND VPWR VPWR tag_array.tag0\[11\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_117_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11507_ clknet_leaf_195_clk _00315_ VGND VGND VPWR VPWR tag_array.tag1\[9\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_152_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12487_ clknet_leaf_240_clk _01181_ VGND VGND VPWR VPWR data_array.data1\[9\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_171_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold109 data_array.data1\[8\]\[14\] VGND VGND VPWR VPWR net1760 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_176_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14226_ clknet_leaf_119_clk _02855_ VGND VGND VPWR VPWR data_array.data1\[12\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_11438_ clknet_leaf_238_clk _00248_ VGND VGND VPWR VPWR data_array.data0\[0\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_153_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_246_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_246_clk
+ sky130_fd_sc_hd__clkbuf_8
X_14157_ clknet_leaf_209_clk _02786_ VGND VGND VPWR VPWR data_array.data0\[2\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_98_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11369_ net1646 net4136 net616 VGND VGND VPWR VPWR _03112_ sky130_fd_sc_hd__mux2_1
XFILLER_4_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_130_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13108_ clknet_leaf_41_clk _01802_ VGND VGND VPWR VPWR data_array.data1\[13\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
X_14088_ clknet_leaf_230_clk _02717_ VGND VGND VPWR VPWR data_array.data0\[1\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_05930_ data_array.rdata0\[33\] net1666 net1147 VGND VGND VPWR VPWR _03414_ sky130_fd_sc_hd__o21a_1
XFILLER_39_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13039_ clknet_leaf_221_clk _01733_ VGND VGND VPWR VPWR data_array.data0\[3\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_85_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1160 net262 VGND VGND VPWR VPWR net1160 sky130_fd_sc_hd__buf_2
XFILLER_152_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1171 net1174 VGND VGND VPWR VPWR net1171 sky130_fd_sc_hd__buf_4
X_05861_ data_array.rdata0\[10\] net852 net1149 VGND VGND VPWR VPWR _03368_ sky130_fd_sc_hd__o21a_1
XFILLER_94_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1182 net1187 VGND VGND VPWR VPWR net1182 sky130_fd_sc_hd__buf_4
Xfanout1193 net1194 VGND VGND VPWR VPWR net1193 sky130_fd_sc_hd__buf_4
X_07600_ data_array.data1\[12\]\[14\] net1381 net1287 data_array.data1\[15\]\[14\]
+ _04826_ VGND VGND VPWR VPWR _04827_ sky130_fd_sc_hd__a221o_1
XFILLER_82_826 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08580_ _03507_ _03509_ net821 VGND VGND VPWR VPWR _05605_ sky130_fd_sc_hd__or3_1
XFILLER_82_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05792_ net2 _03137_ _03252_ _03261_ _03308_ VGND VGND VPWR VPWR _03309_ sky130_fd_sc_hd__a2111o_1
XFILLER_19_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07531_ data_array.data1\[5\]\[8\] net1535 net1439 data_array.data1\[6\]\[8\] VGND
+ VGND VPWR VPWR _04764_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_176_3736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_176_3747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07462_ _04700_ _04701_ VGND VGND VPWR VPWR _00075_ sky130_fd_sc_hd__or2_1
XFILLER_23_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09201_ net777 net4120 net630 VGND VGND VPWR VPWR _00955_ sky130_fd_sc_hd__mux2_1
X_06413_ tag_array.tag0\[1\]\[20\] net1558 net1462 tag_array.tag0\[2\]\[20\] VGND
+ VGND VPWR VPWR _03748_ sky130_fd_sc_hd__a22o_1
X_07393_ data_array.data0\[4\]\[59\] net1379 net1285 data_array.data0\[7\]\[59\] _04638_
+ VGND VGND VPWR VPWR _04639_ sky130_fd_sc_hd__a221o_1
X_09132_ net1014 net3427 net573 VGND VGND VPWR VPWR _00886_ sky130_fd_sc_hd__mux2_1
X_06344_ tag_array.tag0\[4\]\[14\] net1369 net1275 tag_array.tag0\[7\]\[14\] _03684_
+ VGND VGND VPWR VPWR _03685_ sky130_fd_sc_hd__a221o_1
XFILLER_148_677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09063_ net1032 net4279 net414 VGND VGND VPWR VPWR _00817_ sky130_fd_sc_hd__mux2_1
XFILLER_147_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06275_ tag_array.tag0\[9\]\[8\] net1608 net1512 tag_array.tag0\[10\]\[8\] VGND VGND
+ VPWR VPWR _03622_ sky130_fd_sc_hd__a22o_1
XFILLER_148_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08014_ data_array.data1\[12\]\[52\] net1354 net1260 data_array.data1\[15\]\[52\]
+ _05202_ VGND VGND VPWR VPWR _05203_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_7_Left_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold610 data_array.data0\[15\]\[62\] VGND VGND VPWR VPWR net2261 sky130_fd_sc_hd__dlygate4sd3_1
Xhold621 tag_array.tag1\[1\]\[20\] VGND VGND VPWR VPWR net2272 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold632 tag_array.tag1\[11\]\[22\] VGND VGND VPWR VPWR net2283 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_237_clk clknet_5_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_237_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold643 data_array.data1\[8\]\[47\] VGND VGND VPWR VPWR net2294 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold654 tag_array.tag0\[10\]\[21\] VGND VGND VPWR VPWR net2305 sky130_fd_sc_hd__dlygate4sd3_1
Xhold665 tag_array.tag1\[7\]\[19\] VGND VGND VPWR VPWR net2316 sky130_fd_sc_hd__dlygate4sd3_1
Xhold676 data_array.data0\[8\]\[59\] VGND VGND VPWR VPWR net2327 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold687 data_array.data0\[7\]\[7\] VGND VGND VPWR VPWR net2338 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold698 tag_array.tag0\[0\]\[22\] VGND VGND VPWR VPWR net2349 sky130_fd_sc_hd__dlygate4sd3_1
X_09965_ net971 net3743 net370 VGND VGND VPWR VPWR _01714_ sky130_fd_sc_hd__mux2_1
XFILLER_103_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2000 tag_array.tag0\[7\]\[1\] VGND VGND VPWR VPWR net3651 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2011 data_array.data0\[2\]\[57\] VGND VGND VPWR VPWR net3662 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_98_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2022 data_array.data1\[9\]\[41\] VGND VGND VPWR VPWR net3673 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_98_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08916_ net1102 net3002 net428 VGND VGND VPWR VPWR _00672_ sky130_fd_sc_hd__mux2_1
Xhold2033 data_array.data0\[10\]\[8\] VGND VGND VPWR VPWR net3684 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2044 tag_array.tag1\[11\]\[7\] VGND VGND VPWR VPWR net3695 sky130_fd_sc_hd__dlygate4sd3_1
X_09896_ net885 net4075 net379 VGND VGND VPWR VPWR _01646_ sky130_fd_sc_hd__mux2_1
XFILLER_97_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1310 tag_array.tag0\[10\]\[22\] VGND VGND VPWR VPWR net2961 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2055 tag_array.tag0\[0\]\[17\] VGND VGND VPWR VPWR net3706 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2066 data_array.data1\[12\]\[53\] VGND VGND VPWR VPWR net3717 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1321 data_array.data0\[5\]\[59\] VGND VGND VPWR VPWR net2972 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1332 data_array.data1\[14\]\[37\] VGND VGND VPWR VPWR net2983 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2077 data_array.data0\[5\]\[29\] VGND VGND VPWR VPWR net3728 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2088 data_array.data1\[12\]\[20\] VGND VGND VPWR VPWR net3739 sky130_fd_sc_hd__dlygate4sd3_1
X_08847_ net2052 net856 net444 VGND VGND VPWR VPWR _00605_ sky130_fd_sc_hd__mux2_1
Xhold1343 data_array.data0\[3\]\[48\] VGND VGND VPWR VPWR net2994 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1354 data_array.data1\[11\]\[57\] VGND VGND VPWR VPWR net3005 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2099 tag_array.tag0\[6\]\[11\] VGND VGND VPWR VPWR net3750 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1365 data_array.data0\[9\]\[33\] VGND VGND VPWR VPWR net3016 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1376 data_array.data1\[2\]\[8\] VGND VGND VPWR VPWR net3027 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1387 data_array.data1\[15\]\[52\] VGND VGND VPWR VPWR net3038 sky130_fd_sc_hd__dlygate4sd3_1
X_08778_ net712 net3318 net450 VGND VGND VPWR VPWR _00537_ sky130_fd_sc_hd__mux2_1
XFILLER_85_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1398 data_array.data1\[7\]\[24\] VGND VGND VPWR VPWR net3049 sky130_fd_sc_hd__dlygate4sd3_1
X_07729_ data_array.data1\[5\]\[26\] net1525 net1429 data_array.data1\[6\]\[26\] VGND
+ VGND VPWR VPWR _04944_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10740_ net1015 net4322 net499 VGND VGND VPWR VPWR _02485_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10671_ net1731 net1034 net484 VGND VGND VPWR VPWR _02416_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12410_ clknet_leaf_33_clk _01104_ VGND VGND VPWR VPWR data_array.data0\[14\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_13390_ clknet_leaf_118_clk _02020_ VGND VGND VPWR VPWR data_array.data1\[8\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_167_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12341_ clknet_leaf_201_clk _00015_ VGND VGND VPWR VPWR data_array.rdata0\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_182_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12272_ clknet_leaf_194_clk _01030_ VGND VGND VPWR VPWR tag_array.tag1\[13\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_75_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14011_ clknet_leaf_4_clk _02640_ VGND VGND VPWR VPWR data_array.data1\[5\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
X_11223_ net882 net3005 net651 VGND VGND VPWR VPWR _02966_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_228_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_228_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_175_1051 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11154_ net901 net4083 net545 VGND VGND VPWR VPWR _02897_ sky130_fd_sc_hd__mux2_1
XFILLER_136_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10105_ net1765 net702 net638 VGND VGND VPWR VPWR _01854_ sky130_fd_sc_hd__mux2_1
X_11085_ net2244 net920 net334 VGND VGND VPWR VPWR _02828_ sky130_fd_sc_hd__mux2_1
XFILLER_0_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10036_ net942 net3612 net562 VGND VGND VPWR VPWR _01785_ sky130_fd_sc_hd__mux2_1
XFILLER_76_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11987_ clknet_leaf_207_clk _00795_ VGND VGND VPWR VPWR data_array.data0\[4\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13726_ clknet_leaf_24_clk _02355_ VGND VGND VPWR VPWR data_array.data1\[1\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_10938_ net990 net3604 net532 VGND VGND VPWR VPWR _02683_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_154_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_778 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13657_ clknet_leaf_250_clk _02286_ VGND VGND VPWR VPWR data_array.data1\[15\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_10869_ net1008 net2432 net514 VGND VGND VPWR VPWR _02614_ sky130_fd_sc_hd__mux2_1
X_12608_ clknet_leaf_164_clk _01302_ VGND VGND VPWR VPWR tag_array.tag0\[0\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_171_3644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_171_3655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13588_ clknet_leaf_206_clk _02217_ VGND VGND VPWR VPWR data_array.data0\[9\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_30_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12539_ clknet_leaf_101_clk _01233_ VGND VGND VPWR VPWR tag_array.tag1\[11\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_132_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06060_ fsm.tag_out0\[12\] net1120 _03493_ VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__a21o_1
XFILLER_172_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_219_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_219_clk
+ sky130_fd_sc_hd__clkbuf_8
X_14209_ clknet_leaf_234_clk _02838_ VGND VGND VPWR VPWR data_array.data0\[2\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_1018 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout408 net409 VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__clkbuf_8
Xfanout419 net425 VGND VGND VPWR VPWR net419 sky130_fd_sc_hd__clkbuf_4
X_06962_ data_array.data0\[8\]\[20\] net1415 net1321 data_array.data0\[11\]\[20\]
+ _04246_ VGND VGND VPWR VPWR _04247_ sky130_fd_sc_hd__a221o_1
X_09750_ net1844 net787 net667 VGND VGND VPWR VPWR _01502_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05913_ data_array.rdata1\[27\] net830 net839 VGND VGND VPWR VPWR _03403_ sky130_fd_sc_hd__a21o_1
X_08701_ net1726 net718 net489 VGND VGND VPWR VPWR _00460_ sky130_fd_sc_hd__mux2_1
XFILLER_95_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09681_ net763 net3753 net607 VGND VGND VPWR VPWR _01433_ sky130_fd_sc_hd__mux2_1
X_06893_ data_array.data0\[5\]\[14\] net1570 net1474 data_array.data0\[6\]\[14\] VGND
+ VGND VPWR VPWR _04184_ sky130_fd_sc_hd__a22o_1
X_08632_ net694 net4495 net517 VGND VGND VPWR VPWR _00391_ sky130_fd_sc_hd__mux2_1
X_05844_ data_array.rdata1\[4\] net832 net841 VGND VGND VPWR VPWR _03357_ sky130_fd_sc_hd__a21o_1
XFILLER_66_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08563_ net702 net2548 net583 VGND VGND VPWR VPWR _00331_ sky130_fd_sc_hd__mux2_1
XFILLER_54_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05775_ net9 fsm.tag_out1\[10\] VGND VGND VPWR VPWR _03292_ sky130_fd_sc_hd__or2_1
XFILLER_35_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07514_ data_array.data1\[4\]\[6\] net1329 net1235 data_array.data1\[7\]\[6\] _04748_
+ VGND VGND VPWR VPWR _04749_ sky130_fd_sc_hd__a221o_1
XFILLER_35_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08494_ _03507_ _03511_ net822 VGND VGND VPWR VPWR _05566_ sky130_fd_sc_hd__or3_1
XFILLER_22_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07445_ data_array.data1\[9\]\[0\] net1556 net1460 data_array.data1\[10\]\[0\] VGND
+ VGND VPWR VPWR _04686_ sky130_fd_sc_hd__a22o_1
XFILLER_23_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07376_ data_array.data0\[8\]\[58\] net1357 net1263 data_array.data0\[11\]\[58\]
+ _04622_ VGND VGND VPWR VPWR _04623_ sky130_fd_sc_hd__a221o_1
XFILLER_149_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09115_ net1082 net4127 net574 VGND VGND VPWR VPWR _00869_ sky130_fd_sc_hd__mux2_1
XFILLER_13_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06327_ net1637 _03663_ _03667_ net1211 VGND VGND VPWR VPWR _03670_ sky130_fd_sc_hd__a22o_1
XFILLER_109_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09046_ net1102 net2193 net412 VGND VGND VPWR VPWR _00800_ sky130_fd_sc_hd__mux2_1
XFILLER_163_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06258_ tag_array.tag0\[8\]\[6\] net1373 net1279 tag_array.tag0\[11\]\[6\] _03606_
+ VGND VGND VPWR VPWR _03607_ sky130_fd_sc_hd__a221o_1
XFILLER_164_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold440 data_array.data1\[8\]\[29\] VGND VGND VPWR VPWR net2091 sky130_fd_sc_hd__dlygate4sd3_1
X_06189_ tag_array.tag0\[5\]\[0\] net1596 net1500 tag_array.tag0\[6\]\[0\] VGND VGND
+ VPWR VPWR _03544_ sky130_fd_sc_hd__a22o_1
Xhold451 data_array.data0\[0\]\[18\] VGND VGND VPWR VPWR net2102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 data_array.data0\[1\]\[44\] VGND VGND VPWR VPWR net2113 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold473 tag_array.tag0\[4\]\[23\] VGND VGND VPWR VPWR net2124 sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 tag_array.tag1\[0\]\[13\] VGND VGND VPWR VPWR net2135 sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 data_array.data0\[0\]\[40\] VGND VGND VPWR VPWR net2146 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout920 net921 VGND VGND VPWR VPWR net920 sky130_fd_sc_hd__clkbuf_2
Xfanout931 _05510_ VGND VGND VPWR VPWR net931 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_70_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout942 _05504_ VGND VGND VPWR VPWR net942 sky130_fd_sc_hd__clkbuf_2
X_09948_ net1036 net4453 net371 VGND VGND VPWR VPWR _01697_ sky130_fd_sc_hd__mux2_1
Xfanout953 _05498_ VGND VGND VPWR VPWR net953 sky130_fd_sc_hd__buf_1
Xfanout964 net967 VGND VGND VPWR VPWR net964 sky130_fd_sc_hd__clkbuf_2
Xfanout975 _05488_ VGND VGND VPWR VPWR net975 sky130_fd_sc_hd__clkbuf_1
Xfanout986 _05482_ VGND VGND VPWR VPWR net986 sky130_fd_sc_hd__clkbuf_2
X_09879_ net954 net3172 net381 VGND VGND VPWR VPWR _01629_ sky130_fd_sc_hd__mux2_1
Xfanout997 net999 VGND VGND VPWR VPWR net997 sky130_fd_sc_hd__clkbuf_2
Xhold1140 data_array.data1\[5\]\[63\] VGND VGND VPWR VPWR net2791 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1151 data_array.data0\[10\]\[37\] VGND VGND VPWR VPWR net2802 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1162 data_array.data0\[13\]\[62\] VGND VGND VPWR VPWR net2813 sky130_fd_sc_hd__dlygate4sd3_1
X_11910_ clknet_leaf_40_clk _00718_ VGND VGND VPWR VPWR data_array.data0\[5\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1173 data_array.data1\[8\]\[6\] VGND VGND VPWR VPWR net2824 sky130_fd_sc_hd__dlygate4sd3_1
X_12890_ clknet_leaf_207_clk _01584_ VGND VGND VPWR VPWR data_array.data0\[12\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_173_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1184 data_array.data0\[5\]\[56\] VGND VGND VPWR VPWR net2835 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1195 tag_array.tag0\[3\]\[1\] VGND VGND VPWR VPWR net2846 sky130_fd_sc_hd__dlygate4sd3_1
X_11841_ clknet_leaf_47_clk _00649_ VGND VGND VPWR VPWR data_array.data0\[7\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ clknet_leaf_88_clk _00580_ VGND VGND VPWR VPWR data_array.data0\[8\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_68_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10723_ net1083 net4143 net497 VGND VGND VPWR VPWR _02468_ sky130_fd_sc_hd__mux2_1
XFILLER_41_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13511_ clknet_leaf_19_clk _02140_ VGND VGND VPWR VPWR data_array.data1\[0\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_14491_ clknet_leaf_161_clk _03114_ VGND VGND VPWR VPWR tag_array.dirty0\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_9_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13442_ clknet_leaf_121_clk _02072_ VGND VGND VPWR VPWR data_array.data1\[8\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
X_10654_ net1780 net1100 net480 VGND VGND VPWR VPWR _02399_ sky130_fd_sc_hd__mux2_1
XFILLER_167_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13373_ clknet_leaf_180_clk _02003_ VGND VGND VPWR VPWR tag_array.tag0\[2\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_155_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10585_ net864 net3799 net457 VGND VGND VPWR VPWR _02330_ sky130_fd_sc_hd__mux2_1
Xclkload18 clknet_leaf_3_clk VGND VGND VPWR VPWR clkload18/Y sky130_fd_sc_hd__bufinv_16
Xclkload29 clknet_leaf_9_clk VGND VGND VPWR VPWR clkload29/Y sky130_fd_sc_hd__inv_8
XFILLER_103_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12324_ clknet_leaf_269_clk _00060_ VGND VGND VPWR VPWR data_array.rdata0\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_115_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12255_ clknet_leaf_168_clk _01013_ VGND VGND VPWR VPWR tag_array.tag1\[14\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11206_ net951 net3384 net658 VGND VGND VPWR VPWR _02949_ sky130_fd_sc_hd__mux2_1
XFILLER_107_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12186_ clknet_leaf_181_clk _00994_ VGND VGND VPWR VPWR tag_array.tag0\[14\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_122_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11137_ net969 net3245 net541 VGND VGND VPWR VPWR _02880_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_79_Left_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_147_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11068_ net3658 net988 net333 VGND VGND VPWR VPWR _02811_ sky130_fd_sc_hd__mux2_1
XFILLER_62_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10019_ net1010 net2703 net554 VGND VGND VPWR VPWR _01768_ sky130_fd_sc_hd__mux2_1
XFILLER_64_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13709_ clknet_leaf_198_clk _02338_ VGND VGND VPWR VPWR data_array.data1\[1\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_88_Left_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07230_ net1227 _04485_ _04489_ net1179 VGND VGND VPWR VPWR _04491_ sky130_fd_sc_hd__a22o_1
XFILLER_32_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07161_ data_array.data0\[5\]\[38\] net1585 net1489 data_array.data0\[6\]\[38\] VGND
+ VGND VPWR VPWR _04428_ sky130_fd_sc_hd__a22o_1
XFILLER_30_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06112_ data_array.rdata0\[27\] net1136 net1117 data_array.rdata1\[27\] VGND VGND
+ VPWR VPWR net282 sky130_fd_sc_hd__a22o_1
X_07092_ data_array.data0\[0\]\[32\] net1336 net1242 data_array.data0\[3\]\[32\] _04364_
+ VGND VGND VPWR VPWR _04365_ sky130_fd_sc_hd__a221o_1
XFILLER_118_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06043_ net1159 net3 fsm.tag_out1\[4\] net1131 VGND VGND VPWR VPWR _03485_ sky130_fd_sc_hd__a22o_1
XFILLER_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_97_Left_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09802_ net1002 net4036 net389 VGND VGND VPWR VPWR _01553_ sky130_fd_sc_hd__mux2_1
XFILLER_86_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07994_ data_array.data1\[4\]\[50\] net1337 net1243 data_array.data1\[7\]\[50\] _05184_
+ VGND VGND VPWR VPWR _05185_ sky130_fd_sc_hd__a221o_1
X_09733_ net757 net3758 net683 VGND VGND VPWR VPWR _01485_ sky130_fd_sc_hd__mux2_1
X_06945_ _04230_ _04231_ VGND VGND VPWR VPWR _00009_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_2_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09664_ net732 net3734 net613 VGND VGND VPWR VPWR _01416_ sky130_fd_sc_hd__mux2_1
X_06876_ data_array.data0\[4\]\[12\] net1386 net1292 data_array.data0\[7\]\[12\] _04168_
+ VGND VGND VPWR VPWR _04169_ sky130_fd_sc_hd__a221o_1
X_08615_ net764 net3231 net524 VGND VGND VPWR VPWR _00374_ sky130_fd_sc_hd__mux2_1
XFILLER_55_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05827_ _03249_ _03250_ _03259_ _03264_ VGND VGND VPWR VPWR _03344_ sky130_fd_sc_hd__or4_1
X_09595_ net970 net2490 net395 VGND VGND VPWR VPWR _01347_ sky130_fd_sc_hd__mux2_1
XFILLER_83_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08546_ net772 net2990 net588 VGND VGND VPWR VPWR _00314_ sky130_fd_sc_hd__mux2_1
XFILLER_42_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05758_ _03271_ _03272_ _03273_ _03274_ VGND VGND VPWR VPWR _03275_ sky130_fd_sc_hd__or4_1
XFILLER_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1012 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08477_ net824 net813 _05552_ net854 VGND VGND VPWR VPWR _05555_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_46_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05689_ _03203_ _03204_ _03205_ VGND VGND VPWR VPWR _03206_ sky130_fd_sc_hd__or3_1
XFILLER_11_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07428_ net1186 _04665_ _04669_ net1233 VGND VGND VPWR VPWR _04671_ sky130_fd_sc_hd__a22o_1
XFILLER_10_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07359_ data_array.data0\[1\]\[56\] net1533 net1437 data_array.data0\[2\]\[56\] VGND
+ VGND VPWR VPWR _04608_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_21_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_149_Right_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10370_ net720 net4313 net538 VGND VGND VPWR VPWR _02117_ sky130_fd_sc_hd__mux2_1
XFILLER_163_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09029_ net2180 net909 net419 VGND VGND VPWR VPWR _00784_ sky130_fd_sc_hd__mux2_1
XFILLER_124_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12040_ clknet_leaf_241_clk _00848_ VGND VGND VPWR VPWR data_array.data0\[6\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold270 tag_array.tag1\[2\]\[13\] VGND VGND VPWR VPWR net1921 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold281 data_array.data0\[0\]\[52\] VGND VGND VPWR VPWR net1932 sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 data_array.data0\[8\]\[55\] VGND VGND VPWR VPWR net1943 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout750 net753 VGND VGND VPWR VPWR net750 sky130_fd_sc_hd__clkbuf_2
XFILLER_172_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout761 _05381_ VGND VGND VPWR VPWR net761 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout772 net773 VGND VGND VPWR VPWR net772 sky130_fd_sc_hd__clkbuf_2
Xfanout783 _05369_ VGND VGND VPWR VPWR net783 sky130_fd_sc_hd__buf_1
X_13991_ clknet_leaf_36_clk _02620_ VGND VGND VPWR VPWR data_array.data1\[5\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_93_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout794 _05365_ VGND VGND VPWR VPWR net794 sky130_fd_sc_hd__buf_1
XFILLER_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_20 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12942_ clknet_leaf_23_clk _01636_ VGND VGND VPWR VPWR data_array.data0\[13\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12873_ clknet_leaf_260_clk _01567_ VGND VGND VPWR VPWR data_array.data0\[12\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_61_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ clknet_leaf_247_clk _00632_ VGND VGND VPWR VPWR data_array.data0\[7\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_103_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_83_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ clknet_leaf_228_clk _00563_ VGND VGND VPWR VPWR data_array.data0\[8\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_120_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10706_ net2093 net892 net481 VGND VGND VPWR VPWR _02451_ sky130_fd_sc_hd__mux2_1
XFILLER_147_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14474_ clknet_leaf_201_clk _03097_ VGND VGND VPWR VPWR data_array.data1\[7\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11686_ clknet_leaf_32_clk _00494_ VGND VGND VPWR VPWR tag_array.tag1\[15\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_13425_ clknet_leaf_27_clk _02055_ VGND VGND VPWR VPWR data_array.data1\[8\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
X_10637_ net1993 net914 net472 VGND VGND VPWR VPWR _02382_ sky130_fd_sc_hd__mux2_1
Xclkload107 clknet_leaf_32_clk VGND VGND VPWR VPWR clkload107/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload118 clknet_leaf_74_clk VGND VGND VPWR VPWR clkload118/Y sky130_fd_sc_hd__inv_6
Xclkload129 clknet_leaf_85_clk VGND VGND VPWR VPWR clkload129/Y sky130_fd_sc_hd__clkinv_2
X_10568_ net935 net4295 net462 VGND VGND VPWR VPWR _02313_ sky130_fd_sc_hd__mux2_1
X_13356_ clknet_leaf_166_clk _01986_ VGND VGND VPWR VPWR tag_array.tag0\[2\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_116_Right_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12307_ clknet_leaf_231_clk _01065_ VGND VGND VPWR VPWR tag_array.tag1\[12\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_142_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10499_ net949 net3803 net350 VGND VGND VPWR VPWR _02244_ sky130_fd_sc_hd__mux2_1
X_13287_ clknet_leaf_115_clk _01917_ VGND VGND VPWR VPWR data_array.data0\[11\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_149_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12238_ clknet_leaf_183_clk _00168_ VGND VGND VPWR VPWR fsm.tag_out1\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_166_3543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_166_3554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12169_ clknet_leaf_171_clk _00977_ VGND VGND VPWR VPWR tag_array.tag0\[14\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_110_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1909 data_array.data1\[10\]\[51\] VGND VGND VPWR VPWR net3560 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06730_ tag_array.tag1\[9\]\[24\] net1562 net1466 tag_array.tag1\[10\]\[24\] VGND
+ VGND VPWR VPWR _04036_ sky130_fd_sc_hd__a22o_1
Xinput5 cpu_addr[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_2
XFILLER_36_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06661_ tag_array.tag1\[12\]\[18\] net1372 net1278 tag_array.tag1\[15\]\[18\] _03972_
+ VGND VGND VPWR VPWR _03973_ sky130_fd_sc_hd__a221o_1
XFILLER_149_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08400_ net135 net70 net1642 VGND VGND VPWR VPWR _05503_ sky130_fd_sc_hd__mux2_1
XFILLER_18_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05612_ net1649 VGND VGND VPWR VPWR _03134_ sky130_fd_sc_hd__inv_2
XFILLER_52_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09380_ net880 net4129 net405 VGND VGND VPWR VPWR _01133_ sky130_fd_sc_hd__mux2_1
X_06592_ net1187 _03905_ _03909_ net1234 VGND VGND VPWR VPWR _03911_ sky130_fd_sc_hd__a22o_1
XFILLER_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08331_ net109 net44 net1641 VGND VGND VPWR VPWR _05457_ sky130_fd_sc_hd__mux2_1
XFILLER_33_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08262_ net703 net2876 net798 VGND VGND VPWR VPWR _00218_ sky130_fd_sc_hd__mux2_1
XFILLER_119_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07213_ data_array.data0\[0\]\[43\] net1378 net1284 data_array.data0\[3\]\[43\] _04474_
+ VGND VGND VPWR VPWR _04475_ sky130_fd_sc_hd__a221o_1
X_08193_ net1650 net1161 net30 VGND VGND VPWR VPWR _05363_ sky130_fd_sc_hd__and3_1
XFILLER_119_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07144_ data_array.data0\[9\]\[37\] net1547 net1451 data_array.data0\[10\]\[37\]
+ VGND VGND VPWR VPWR _04412_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_41_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1046 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07075_ net1630 _04343_ _04347_ net1204 VGND VGND VPWR VPWR _04350_ sky130_fd_sc_hd__a22o_1
Xoutput320 net320 VGND VGND VPWR VPWR mem_wdata[61] sky130_fd_sc_hd__buf_2
XFILLER_126_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06026_ fsm.lru_out net327 VGND VGND VPWR VPWR _03476_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_7_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07977_ net1630 _05163_ _05167_ net1204 VGND VGND VPWR VPWR _05170_ sky130_fd_sc_hd__a22o_1
XFILLER_75_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_87_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09716_ net722 net3516 net610 VGND VGND VPWR VPWR _01468_ sky130_fd_sc_hd__mux2_1
X_06928_ data_array.data0\[9\]\[17\] net1528 net1432 data_array.data0\[10\]\[17\]
+ VGND VGND VPWR VPWR _04216_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_87_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09647_ net698 net3576 net616 VGND VGND VPWR VPWR _01399_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06859_ data_array.data0\[8\]\[11\] net1383 net1289 data_array.data0\[11\]\[11\]
+ _04152_ VGND VGND VPWR VPWR _04153_ sky130_fd_sc_hd__a221o_1
XFILLER_43_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09578_ net1037 net3376 net395 VGND VGND VPWR VPWR _01330_ sky130_fd_sc_hd__mux2_1
XFILLER_43_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08529_ net814 _05590_ VGND VGND VPWR VPWR _05591_ sky130_fd_sc_hd__nand2_2
XFILLER_51_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11540_ clknet_leaf_193_clk _00348_ VGND VGND VPWR VPWR tag_array.tag1\[6\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_51_692 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11471_ clknet_leaf_114_clk _00281_ VGND VGND VPWR VPWR data_array.data0\[0\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13210_ clknet_leaf_80_clk _00105_ VGND VGND VPWR VPWR data_array.rdata1\[47\] sky130_fd_sc_hd__dfxtp_1
X_10422_ net2047 net965 net668 VGND VGND VPWR VPWR _02168_ sky130_fd_sc_hd__mux2_1
XFILLER_136_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14190_ clknet_leaf_87_clk _02819_ VGND VGND VPWR VPWR data_array.data0\[2\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13141_ clknet_leaf_191_clk _01835_ VGND VGND VPWR VPWR tag_array.tag1\[8\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_10353_ net790 net4080 net538 VGND VGND VPWR VPWR _02100_ sky130_fd_sc_hd__mux2_1
XFILLER_3_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13072_ clknet_leaf_204_clk _01766_ VGND VGND VPWR VPWR data_array.data1\[13\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_10284_ net2011 net1025 net637 VGND VGND VPWR VPWR _02031_ sky130_fd_sc_hd__mux2_1
XFILLER_140_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12023_ clknet_leaf_90_clk _00831_ VGND VGND VPWR VPWR data_array.data0\[6\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout1501 net1504 VGND VGND VPWR VPWR net1501 sky130_fd_sc_hd__clkbuf_4
Xfanout1512 net1513 VGND VGND VPWR VPWR net1512 sky130_fd_sc_hd__clkbuf_4
Xfanout1523 net1524 VGND VGND VPWR VPWR net1523 sky130_fd_sc_hd__clkbuf_4
XFILLER_132_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1534 net1536 VGND VGND VPWR VPWR net1534 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_144_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1545 net1546 VGND VGND VPWR VPWR net1545 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_144_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1556 net1557 VGND VGND VPWR VPWR net1556 sky130_fd_sc_hd__clkbuf_4
XFILLER_78_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1567 net1569 VGND VGND VPWR VPWR net1567 sky130_fd_sc_hd__clkbuf_4
Xfanout580 net581 VGND VGND VPWR VPWR net580 sky130_fd_sc_hd__clkbuf_8
Xfanout1578 net1579 VGND VGND VPWR VPWR net1578 sky130_fd_sc_hd__clkbuf_2
Xfanout1589 net1590 VGND VGND VPWR VPWR net1589 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_161_3451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout591 net594 VGND VGND VPWR VPWR net591 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_161_3462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13974_ clknet_leaf_51_clk _02603_ VGND VGND VPWR VPWR data_array.data1\[5\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_122_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12925_ clknet_leaf_55_clk _01619_ VGND VGND VPWR VPWR data_array.data0\[13\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12856_ clknet_leaf_97_clk _01550_ VGND VGND VPWR VPWR data_array.data0\[12\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_11807_ clknet_leaf_61_clk _00615_ VGND VGND VPWR VPWR data_array.data0\[7\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12787_ clknet_leaf_134_clk _01481_ VGND VGND VPWR VPWR tag_array.tag1\[10\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_159_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11738_ clknet_leaf_73_clk _00546_ VGND VGND VPWR VPWR data_array.data0\[8\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_147_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_848 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14457_ clknet_leaf_258_clk _03080_ VGND VGND VPWR VPWR data_array.data1\[7\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
X_11669_ clknet_leaf_102_clk _00477_ VGND VGND VPWR VPWR tag_array.tag1\[1\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_13408_ clknet_leaf_30_clk _02038_ VGND VGND VPWR VPWR data_array.data1\[8\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_14388_ clknet_leaf_77_clk _03011_ VGND VGND VPWR VPWR data_array.data1\[10\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_127_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13339_ clknet_leaf_56_clk _01969_ VGND VGND VPWR VPWR data_array.data0\[10\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_182_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07900_ net1616 _05093_ _05097_ net1190 VGND VGND VPWR VPWR _05100_ sky130_fd_sc_hd__a22o_1
XFILLER_29_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2407 data_array.data0\[15\]\[23\] VGND VGND VPWR VPWR net4058 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2418 data_array.data1\[6\]\[4\] VGND VGND VPWR VPWR net4069 sky130_fd_sc_hd__dlygate4sd3_1
X_08880_ net986 net4005 net439 VGND VGND VPWR VPWR _00637_ sky130_fd_sc_hd__mux2_1
XFILLER_29_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_181_3838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2429 tag_array.tag0\[15\]\[1\] VGND VGND VPWR VPWR net4080 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1706 data_array.data1\[8\]\[23\] VGND VGND VPWR VPWR net3357 sky130_fd_sc_hd__dlygate4sd3_1
X_07831_ data_array.data1\[8\]\[35\] net1336 net1242 data_array.data1\[11\]\[35\]
+ _05036_ VGND VGND VPWR VPWR _05037_ sky130_fd_sc_hd__a221o_1
Xhold1717 data_array.data1\[13\]\[41\] VGND VGND VPWR VPWR net3368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1728 data_array.data1\[10\]\[21\] VGND VGND VPWR VPWR net3379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1739 data_array.data1\[7\]\[16\] VGND VGND VPWR VPWR net3390 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07762_ data_array.data1\[1\]\[29\] net1573 net1477 data_array.data1\[2\]\[29\] VGND
+ VGND VPWR VPWR _04974_ sky130_fd_sc_hd__a22o_1
XFILLER_38_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09501_ net723 net3058 net625 VGND VGND VPWR VPWR _01254_ sky130_fd_sc_hd__mux2_1
X_06713_ net1220 _04015_ _04019_ net1171 VGND VGND VPWR VPWR _04021_ sky130_fd_sc_hd__a22o_1
X_07693_ _04910_ _04911_ VGND VGND VPWR VPWR _00078_ sky130_fd_sc_hd__or2_1
XFILLER_65_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06644_ tag_array.tag1\[5\]\[16\] net1609 net1513 tag_array.tag1\[6\]\[16\] VGND
+ VGND VPWR VPWR _03958_ sky130_fd_sc_hd__a22o_1
X_09432_ net937 net3249 net585 VGND VGND VPWR VPWR _01185_ sky130_fd_sc_hd__mux2_1
XFILLER_52_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09363_ net948 net2202 net408 VGND VGND VPWR VPWR _01116_ sky130_fd_sc_hd__mux2_1
X_06575_ tag_array.tag1\[0\]\[10\] net1404 net1310 tag_array.tag1\[3\]\[10\] _03894_
+ VGND VGND VPWR VPWR _03895_ sky130_fd_sc_hd__a221o_1
XFILLER_178_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08314_ net1126 _05445_ VGND VGND VPWR VPWR _05446_ sky130_fd_sc_hd__and2_2
X_09294_ net703 net3130 net558 VGND VGND VPWR VPWR _01048_ sky130_fd_sc_hd__mux2_1
XANTENNA_10 _00158_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 _03506_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_32 net334 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08245_ net1651 net1163 net17 VGND VGND VPWR VPWR _05398_ sky130_fd_sc_hd__and3_1
XANTENNA_43 net532 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_54 net1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_65 net1624 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_76 net369 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_87 net1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08176_ net1174 _05345_ _05349_ net1223 VGND VGND VPWR VPWR _05351_ sky130_fd_sc_hd__a22o_1
XFILLER_119_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07127_ data_array.data0\[8\]\[35\] net1346 net1252 data_array.data0\[11\]\[35\]
+ _04396_ VGND VGND VPWR VPWR _04397_ sky130_fd_sc_hd__a221o_1
XFILLER_173_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07058_ data_array.data0\[1\]\[29\] net1571 net1475 data_array.data0\[2\]\[29\] VGND
+ VGND VPWR VPWR _04334_ sky130_fd_sc_hd__a22o_1
XFILLER_161_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput172 net172 VGND VGND VPWR VPWR cpu_rdata[16] sky130_fd_sc_hd__clkbuf_4
X_06009_ data_array.rdata1\[59\] net833 net842 VGND VGND VPWR VPWR _03467_ sky130_fd_sc_hd__a21o_1
Xoutput183 net183 VGND VGND VPWR VPWR cpu_rdata[26] sky130_fd_sc_hd__buf_4
XFILLER_82_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput194 net194 VGND VGND VPWR VPWR cpu_rdata[36] sky130_fd_sc_hd__buf_2
XFILLER_43_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2930 tag_array.tag1\[9\]\[6\] VGND VGND VPWR VPWR net4581 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2941 data_array.data1\[10\]\[57\] VGND VGND VPWR VPWR net4592 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_153_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2952 data_array.data0\[12\]\[28\] VGND VGND VPWR VPWR net4603 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2963 fsm.state\[3\] VGND VGND VPWR VPWR net4614 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2974 fsm.state\[5\] VGND VGND VPWR VPWR net4625 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_16_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10971_ net858 net3708 net528 VGND VGND VPWR VPWR _02716_ sky130_fd_sc_hd__mux2_1
XFILLER_29_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12710_ clknet_leaf_178_clk _01404_ VGND VGND VPWR VPWR tag_array.tag0\[7\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_13690_ clknet_leaf_245_clk _02319_ VGND VGND VPWR VPWR data_array.data1\[15\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_71_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12641_ clknet_leaf_176_clk _01335_ VGND VGND VPWR VPWR data_array.data0\[15\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12572_ clknet_leaf_178_clk _01266_ VGND VGND VPWR VPWR tag_array.tag0\[10\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_178_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14311_ clknet_leaf_37_clk _02940_ VGND VGND VPWR VPWR data_array.data1\[11\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_11523_ clknet_leaf_197_clk _00331_ VGND VGND VPWR VPWR tag_array.tag1\[9\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14242_ clknet_leaf_255_clk _02871_ VGND VGND VPWR VPWR data_array.data1\[12\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_11454_ clknet_leaf_48_clk _00264_ VGND VGND VPWR VPWR data_array.data0\[0\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_172_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10405_ net1742 net1034 net668 VGND VGND VPWR VPWR _02151_ sky130_fd_sc_hd__mux2_1
XFILLER_183_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14173_ clknet_leaf_226_clk _02802_ VGND VGND VPWR VPWR data_array.data0\[2\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_11385_ clknet_leaf_175_clk _00195_ VGND VGND VPWR VPWR lru_array.lru_mem\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_152_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13124_ clknet_leaf_165_clk _01818_ VGND VGND VPWR VPWR tag_array.tag0\[3\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_10336_ net754 net4417 net593 VGND VGND VPWR VPWR _02083_ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_9_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_9_0_clk sky130_fd_sc_hd__clkbuf_8
X_10267_ net2391 net1094 net640 VGND VGND VPWR VPWR _02014_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_163_3502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13055_ clknet_leaf_268_clk _01749_ VGND VGND VPWR VPWR data_array.data1\[13\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1320 net1322 VGND VGND VPWR VPWR net1320 sky130_fd_sc_hd__clkbuf_4
XFILLER_121_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12006_ clknet_leaf_223_clk _00814_ VGND VGND VPWR VPWR data_array.data0\[6\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_39_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1331 net1376 VGND VGND VPWR VPWR net1331 sky130_fd_sc_hd__buf_2
Xfanout1342 net1352 VGND VGND VPWR VPWR net1342 sky130_fd_sc_hd__clkbuf_2
XFILLER_94_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10198_ net1012 net2657 net358 VGND VGND VPWR VPWR _01945_ sky130_fd_sc_hd__mux2_1
XFILLER_120_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1353 net1355 VGND VGND VPWR VPWR net1353 sky130_fd_sc_hd__clkbuf_4
Xfanout1364 net1376 VGND VGND VPWR VPWR net1364 sky130_fd_sc_hd__clkbuf_4
XFILLER_94_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1375 net1376 VGND VGND VPWR VPWR net1375 sky130_fd_sc_hd__clkbuf_2
Xfanout1386 net1387 VGND VGND VPWR VPWR net1386 sky130_fd_sc_hd__clkbuf_4
Xfanout1397 net1398 VGND VGND VPWR VPWR net1397 sky130_fd_sc_hd__clkbuf_4
X_13957_ clknet_leaf_211_clk _02586_ VGND VGND VPWR VPWR data_array.data1\[4\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
X_12908_ clknet_leaf_94_clk _01602_ VGND VGND VPWR VPWR data_array.data0\[13\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13888_ clknet_leaf_8_clk _02517_ VGND VGND VPWR VPWR data_array.data1\[3\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12839_ clknet_leaf_113_clk _01533_ VGND VGND VPWR VPWR data_array.data0\[12\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06360_ net1207 _03693_ _03697_ net1633 VGND VGND VPWR VPWR _03700_ sky130_fd_sc_hd__a22o_1
XFILLER_159_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06291_ tag_array.tag0\[8\]\[9\] net1409 net1315 tag_array.tag0\[11\]\[9\] _03636_
+ VGND VGND VPWR VPWR _03637_ sky130_fd_sc_hd__a221o_1
XFILLER_174_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08030_ data_array.data1\[5\]\[53\] net1524 net1428 data_array.data1\[6\]\[53\] VGND
+ VGND VPWR VPWR _05218_ sky130_fd_sc_hd__a22o_1
Xinput30 cpu_addr[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_135_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput41 cpu_wdata[16] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_135_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput52 cpu_wdata[26] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_1
XFILLER_116_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput63 cpu_wdata[36] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_1
XFILLER_162_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold803 data_array.data0\[13\]\[5\] VGND VGND VPWR VPWR net2454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold814 data_array.data1\[2\]\[37\] VGND VGND VPWR VPWR net2465 sky130_fd_sc_hd__dlygate4sd3_1
Xinput74 cpu_wdata[46] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_1
XFILLER_116_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput85 cpu_wdata[56] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_1
Xhold825 data_array.data1\[1\]\[55\] VGND VGND VPWR VPWR net2476 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput96 cpu_wdata[8] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_1
XFILLER_66_1016 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold836 tag_array.tag0\[9\]\[8\] VGND VGND VPWR VPWR net2487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold847 data_array.data0\[5\]\[36\] VGND VGND VPWR VPWR net2498 sky130_fd_sc_hd__dlygate4sd3_1
Xhold858 data_array.data1\[11\]\[50\] VGND VGND VPWR VPWR net2509 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09981_ net904 net4452 net370 VGND VGND VPWR VPWR _01730_ sky130_fd_sc_hd__mux2_1
XFILLER_104_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold869 data_array.data0\[7\]\[33\] VGND VGND VPWR VPWR net2520 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08932_ net1036 net3128 net431 VGND VGND VPWR VPWR _00688_ sky130_fd_sc_hd__mux2_1
XFILLER_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2204 data_array.data0\[14\]\[58\] VGND VGND VPWR VPWR net3855 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2215 tag_array.tag1\[5\]\[2\] VGND VGND VPWR VPWR net3866 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2226 data_array.data0\[3\]\[7\] VGND VGND VPWR VPWR net3877 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2237 data_array.data1\[2\]\[32\] VGND VGND VPWR VPWR net3888 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_36_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1503 data_array.data0\[10\]\[35\] VGND VGND VPWR VPWR net3154 sky130_fd_sc_hd__dlygate4sd3_1
X_08863_ net1052 net4305 net439 VGND VGND VPWR VPWR _00620_ sky130_fd_sc_hd__mux2_1
Xhold2248 tag_array.tag1\[11\]\[11\] VGND VGND VPWR VPWR net3899 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2259 data_array.data1\[11\]\[44\] VGND VGND VPWR VPWR net3910 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1514 data_array.data1\[13\]\[46\] VGND VGND VPWR VPWR net3165 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1525 data_array.data1\[4\]\[20\] VGND VGND VPWR VPWR net3176 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_24_Left_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07814_ _05020_ _05021_ VGND VGND VPWR VPWR _00090_ sky130_fd_sc_hd__or2_1
Xhold1536 data_array.data1\[14\]\[26\] VGND VGND VPWR VPWR net3187 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1547 data_array.data1\[14\]\[44\] VGND VGND VPWR VPWR net3198 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1558 data_array.data1\[6\]\[8\] VGND VGND VPWR VPWR net3209 sky130_fd_sc_hd__dlygate4sd3_1
X_08794_ net2097 net1069 net448 VGND VGND VPWR VPWR _00552_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_84_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1569 data_array.data1\[9\]\[11\] VGND VGND VPWR VPWR net3220 sky130_fd_sc_hd__dlygate4sd3_1
X_07745_ data_array.data1\[4\]\[27\] net1356 net1262 data_array.data1\[7\]\[27\] _04958_
+ VGND VGND VPWR VPWR _04959_ sky130_fd_sc_hd__a221o_1
XFILLER_65_581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07676_ data_array.data1\[13\]\[21\] net1547 net1451 data_array.data1\[14\]\[21\]
+ VGND VGND VPWR VPWR _04896_ sky130_fd_sc_hd__a22o_1
X_09415_ net1005 net2950 net579 VGND VGND VPWR VPWR _01168_ sky130_fd_sc_hd__mux2_1
XFILLER_41_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06627_ tag_array.tag1\[9\]\[15\] net1592 net1496 tag_array.tag1\[10\]\[15\] VGND
+ VGND VPWR VPWR _03942_ sky130_fd_sc_hd__a22o_1
XFILLER_179_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09346_ net1019 net3994 net404 VGND VGND VPWR VPWR _01099_ sky130_fd_sc_hd__mux2_1
X_06558_ net1636 _03873_ _03877_ net1210 VGND VGND VPWR VPWR _03880_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_33_Left_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09277_ net773 net3144 net564 VGND VGND VPWR VPWR _01031_ sky130_fd_sc_hd__mux2_1
X_06489_ tag_array.tag1\[12\]\[2\] net1349 net1255 tag_array.tag1\[15\]\[2\] _03816_
+ VGND VGND VPWR VPWR _03817_ sky130_fd_sc_hd__a221o_1
XFILLER_166_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08228_ fsm.tag_out1\[11\] net818 net810 fsm.tag_out0\[11\] _05386_ VGND VGND VPWR
+ VPWR _05387_ sky130_fd_sc_hd__a221o_4
XFILLER_165_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08159_ tag_array.dirty0\[0\] net1403 net1309 tag_array.dirty0\[3\] _05334_ VGND
+ VGND VPWR VPWR _05335_ sky130_fd_sc_hd__a221o_1
XFILLER_134_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11170_ net1095 net4124 net656 VGND VGND VPWR VPWR _02913_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10121_ net1060 net2313 net368 VGND VGND VPWR VPWR _01869_ sky130_fd_sc_hd__mux2_1
XFILLER_0_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_42_Left_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10052_ net879 net3362 net558 VGND VGND VPWR VPWR _01801_ sky130_fd_sc_hd__mux2_1
XFILLER_76_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_995 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2760 data_array.data1\[10\]\[30\] VGND VGND VPWR VPWR net4411 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2771 data_array.data0\[13\]\[38\] VGND VGND VPWR VPWR net4422 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2782 data_array.data0\[13\]\[53\] VGND VGND VPWR VPWR net4433 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2793 data_array.data1\[7\]\[46\] VGND VGND VPWR VPWR net4444 sky130_fd_sc_hd__dlygate4sd3_1
X_13811_ clknet_leaf_36_clk _02440_ VGND VGND VPWR VPWR data_array.data1\[2\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_180_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13742_ clknet_leaf_74_clk _02371_ VGND VGND VPWR VPWR data_array.data1\[1\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
X_10954_ net924 net4528 net526 VGND VGND VPWR VPWR _02699_ sky130_fd_sc_hd__mux2_1
XFILLER_73_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13673_ clknet_leaf_75_clk _02302_ VGND VGND VPWR VPWR data_array.data1\[15\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_139_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10885_ net944 net3008 net514 VGND VGND VPWR VPWR _02630_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_191_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_191_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_139_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1040 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Left_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12624_ clknet_leaf_0_clk _01318_ VGND VGND VPWR VPWR data_array.data0\[15\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_169_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12555_ clknet_leaf_153_clk _01249_ VGND VGND VPWR VPWR tag_array.tag0\[11\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_117_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11506_ clknet_leaf_134_clk _00314_ VGND VGND VPWR VPWR tag_array.tag1\[9\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_172_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12486_ clknet_leaf_77_clk _01180_ VGND VGND VPWR VPWR data_array.data1\[9\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
X_14225_ clknet_leaf_57_clk _02854_ VGND VGND VPWR VPWR data_array.data1\[12\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_11437_ clknet_leaf_246_clk _00247_ VGND VGND VPWR VPWR data_array.data0\[0\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_171_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14156_ clknet_leaf_57_clk _02785_ VGND VGND VPWR VPWR data_array.data0\[2\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_11368_ net1646 net3990 net613 VGND VGND VPWR VPWR _03111_ sky130_fd_sc_hd__mux2_1
XFILLER_140_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13107_ clknet_leaf_203_clk _01801_ VGND VGND VPWR VPWR data_array.data1\[13\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_60_Left_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10319_ net2844 net887 net635 VGND VGND VPWR VPWR _02066_ sky130_fd_sc_hd__mux2_1
X_14087_ clknet_leaf_204_clk _02716_ VGND VGND VPWR VPWR data_array.data1\[6\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
X_11299_ net1098 net4448 net800 VGND VGND VPWR VPWR _03042_ sky130_fd_sc_hd__mux2_1
XFILLER_112_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13038_ clknet_leaf_3_clk _01732_ VGND VGND VPWR VPWR data_array.data0\[3\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_79_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1150 net1151 VGND VGND VPWR VPWR net1150 sky130_fd_sc_hd__buf_4
XFILLER_121_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05860_ net162 net1155 _03366_ _03367_ VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__a22o_1
Xfanout1161 net1162 VGND VGND VPWR VPWR net1161 sky130_fd_sc_hd__buf_2
XFILLER_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1172 net1174 VGND VGND VPWR VPWR net1172 sky130_fd_sc_hd__buf_4
Xfanout1183 net1186 VGND VGND VPWR VPWR net1183 sky130_fd_sc_hd__buf_4
Xfanout1194 net1212 VGND VGND VPWR VPWR net1194 sky130_fd_sc_hd__clkbuf_4
XFILLER_81_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05791_ net19 fsm.tag_out1\[19\] VGND VGND VPWR VPWR _03308_ sky130_fd_sc_hd__and2b_1
XFILLER_82_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07530_ data_array.data1\[12\]\[8\] net1344 net1250 data_array.data1\[15\]\[8\] _04762_
+ VGND VGND VPWR VPWR _04763_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_176_3737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07461_ net1213 _04695_ _04699_ net1165 VGND VGND VPWR VPWR _04701_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_176_3748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_182_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_182_clk
+ sky130_fd_sc_hd__clkbuf_8
X_06412_ tag_array.tag0\[8\]\[20\] net1369 net1276 tag_array.tag0\[11\]\[20\] _03746_
+ VGND VGND VPWR VPWR _03747_ sky130_fd_sc_hd__a221o_1
X_09200_ net781 net3116 net630 VGND VGND VPWR VPWR _00954_ sky130_fd_sc_hd__mux2_1
XFILLER_167_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07392_ data_array.data0\[5\]\[59\] net1570 net1474 data_array.data0\[6\]\[59\] VGND
+ VGND VPWR VPWR _04638_ sky130_fd_sc_hd__a22o_1
XFILLER_33_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09131_ net1016 net3549 net570 VGND VGND VPWR VPWR _00885_ sky130_fd_sc_hd__mux2_1
X_06343_ tag_array.tag0\[5\]\[14\] net1559 net1463 tag_array.tag0\[6\]\[14\] VGND
+ VGND VPWR VPWR _03684_ sky130_fd_sc_hd__a22o_1
XFILLER_148_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09062_ net1036 net3342 net415 VGND VGND VPWR VPWR _00816_ sky130_fd_sc_hd__mux2_1
X_06274_ _03620_ _03621_ VGND VGND VPWR VPWR _00153_ sky130_fd_sc_hd__or2_1
XFILLER_148_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08013_ data_array.data1\[13\]\[52\] net1546 net1450 data_array.data1\[14\]\[52\]
+ VGND VGND VPWR VPWR _05202_ sky130_fd_sc_hd__a22o_1
XFILLER_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold600 data_array.data1\[0\]\[27\] VGND VGND VPWR VPWR net2251 sky130_fd_sc_hd__dlygate4sd3_1
Xhold611 data_array.data1\[1\]\[14\] VGND VGND VPWR VPWR net2262 sky130_fd_sc_hd__dlygate4sd3_1
Xhold622 data_array.data0\[0\]\[50\] VGND VGND VPWR VPWR net2273 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold633 tag_array.tag1\[3\]\[18\] VGND VGND VPWR VPWR net2284 sky130_fd_sc_hd__dlygate4sd3_1
Xhold644 data_array.data0\[10\]\[15\] VGND VGND VPWR VPWR net2295 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold655 tag_array.tag1\[4\]\[7\] VGND VGND VPWR VPWR net2306 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold666 data_array.data0\[2\]\[49\] VGND VGND VPWR VPWR net2317 sky130_fd_sc_hd__dlygate4sd3_1
Xhold677 data_array.data0\[4\]\[34\] VGND VGND VPWR VPWR net2328 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold688 tag_array.tag1\[4\]\[20\] VGND VGND VPWR VPWR net2339 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold699 data_array.data1\[2\]\[50\] VGND VGND VPWR VPWR net2350 sky130_fd_sc_hd__dlygate4sd3_1
X_09964_ net972 net4057 net370 VGND VGND VPWR VPWR _01713_ sky130_fd_sc_hd__mux2_1
Xhold2001 data_array.data1\[13\]\[57\] VGND VGND VPWR VPWR net3652 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2012 data_array.data1\[7\]\[62\] VGND VGND VPWR VPWR net3663 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08915_ net1106 net3363 net426 VGND VGND VPWR VPWR _00671_ sky130_fd_sc_hd__mux2_1
Xhold2023 data_array.data1\[5\]\[46\] VGND VGND VPWR VPWR net3674 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2034 data_array.data0\[15\]\[45\] VGND VGND VPWR VPWR net3685 sky130_fd_sc_hd__dlygate4sd3_1
X_09895_ net889 net2736 net379 VGND VGND VPWR VPWR _01645_ sky130_fd_sc_hd__mux2_1
Xhold2045 data_array.data0\[6\]\[58\] VGND VGND VPWR VPWR net3696 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1300 data_array.data0\[15\]\[56\] VGND VGND VPWR VPWR net2951 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1311 data_array.data0\[2\]\[32\] VGND VGND VPWR VPWR net2962 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2056 data_array.data0\[9\]\[7\] VGND VGND VPWR VPWR net3707 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1322 data_array.data0\[12\]\[29\] VGND VGND VPWR VPWR net2973 sky130_fd_sc_hd__dlygate4sd3_1
X_08846_ net1836 net861 net449 VGND VGND VPWR VPWR _00604_ sky130_fd_sc_hd__mux2_1
Xhold2067 data_array.data0\[10\]\[25\] VGND VGND VPWR VPWR net3718 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1333 data_array.data1\[12\]\[4\] VGND VGND VPWR VPWR net2984 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2078 data_array.data1\[12\]\[63\] VGND VGND VPWR VPWR net3729 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1344 data_array.data1\[5\]\[19\] VGND VGND VPWR VPWR net2995 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2089 data_array.data0\[15\]\[63\] VGND VGND VPWR VPWR net3740 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1355 tag_array.tag1\[5\]\[6\] VGND VGND VPWR VPWR net3006 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1366 data_array.data0\[13\]\[61\] VGND VGND VPWR VPWR net3017 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1377 data_array.data0\[2\]\[7\] VGND VGND VPWR VPWR net3028 sky130_fd_sc_hd__dlygate4sd3_1
X_08777_ net717 net4385 net451 VGND VGND VPWR VPWR _00536_ sky130_fd_sc_hd__mux2_1
Xhold1388 data_array.data0\[1\]\[1\] VGND VGND VPWR VPWR net3039 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_05989_ net146 net1152 _03452_ _03453_ VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_108_Left_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1399 data_array.data0\[10\]\[9\] VGND VGND VPWR VPWR net3050 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07728_ data_array.data1\[8\]\[26\] net1335 net1241 data_array.data1\[11\]\[26\]
+ _04942_ VGND VGND VPWR VPWR _04943_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_0_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07659_ net1178 _04875_ _04879_ net1226 VGND VGND VPWR VPWR _04881_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_173_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_173_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_81_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10670_ net2088 net1038 net483 VGND VGND VPWR VPWR _02415_ sky130_fd_sc_hd__mux2_1
X_09329_ net1084 net4325 net402 VGND VGND VPWR VPWR _01082_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12340_ clknet_leaf_12_clk _00014_ VGND VGND VPWR VPWR data_array.rdata0\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12271_ clknet_leaf_191_clk _01029_ VGND VGND VPWR VPWR tag_array.tag1\[13\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_182_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14010_ clknet_leaf_245_clk _02639_ VGND VGND VPWR VPWR data_array.data1\[5\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_75_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11222_ net887 net2710 net650 VGND VGND VPWR VPWR _02965_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_112_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11153_ net907 net3181 net541 VGND VGND VPWR VPWR _02896_ sky130_fd_sc_hd__mux2_1
XFILLER_122_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10104_ net2017 net707 net643 VGND VGND VPWR VPWR _01853_ sky130_fd_sc_hd__mux2_1
X_11084_ net2105 net926 net328 VGND VGND VPWR VPWR _02827_ sky130_fd_sc_hd__mux2_1
XFILLER_0_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10035_ net947 net3368 net554 VGND VGND VPWR VPWR _01784_ sky130_fd_sc_hd__mux2_1
XFILLER_76_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2590 data_array.data1\[5\]\[51\] VGND VGND VPWR VPWR net4241 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11986_ clknet_leaf_110_clk _00794_ VGND VGND VPWR VPWR data_array.data0\[4\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13725_ clknet_leaf_228_clk _02354_ VGND VGND VPWR VPWR data_array.data1\[1\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_10937_ net994 net2759 net531 VGND VGND VPWR VPWR _02682_ sky130_fd_sc_hd__mux2_1
XFILLER_56_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_164_clk clknet_5_25__leaf_clk VGND VGND VPWR VPWR clknet_leaf_164_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_44_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13656_ clknet_leaf_213_clk _02285_ VGND VGND VPWR VPWR data_array.data1\[15\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10868_ net1014 net3019 net520 VGND VGND VPWR VPWR _02613_ sky130_fd_sc_hd__mux2_1
X_12607_ clknet_leaf_169_clk _01301_ VGND VGND VPWR VPWR tag_array.tag0\[0\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_129_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13587_ clknet_leaf_94_clk _02216_ VGND VGND VPWR VPWR data_array.data0\[9\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_171_3656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10799_ net1818 net1034 net508 VGND VGND VPWR VPWR _02544_ sky130_fd_sc_hd__mux2_1
XFILLER_158_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12538_ clknet_leaf_232_clk _01232_ VGND VGND VPWR VPWR tag_array.tag1\[11\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_118_829 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1070 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12469_ clknet_leaf_221_clk _01163_ VGND VGND VPWR VPWR data_array.data1\[9\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_173_979 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14208_ clknet_leaf_12_clk _02837_ VGND VGND VPWR VPWR data_array.data0\[2\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14139_ clknet_leaf_2_clk _02768_ VGND VGND VPWR VPWR data_array.data0\[1\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout409 _03123_ VGND VGND VPWR VPWR net409 sky130_fd_sc_hd__buf_4
X_06961_ data_array.data0\[9\]\[20\] net1605 net1509 data_array.data0\[10\]\[20\]
+ VGND VGND VPWR VPWR _04246_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_33_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08700_ net2132 net724 net487 VGND VGND VPWR VPWR _00459_ sky130_fd_sc_hd__mux2_1
X_05912_ data_array.rdata0\[27\] net848 net1144 VGND VGND VPWR VPWR _03402_ sky130_fd_sc_hd__o21a_1
X_09680_ net768 net4257 net605 VGND VGND VPWR VPWR _01432_ sky130_fd_sc_hd__mux2_1
XFILLER_104_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06892_ data_array.data0\[8\]\[14\] net1378 net1284 data_array.data0\[11\]\[14\]
+ _04182_ VGND VGND VPWR VPWR _04183_ sky130_fd_sc_hd__a221o_1
XFILLER_95_985 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08631_ net700 net4072 net524 VGND VGND VPWR VPWR _00390_ sky130_fd_sc_hd__mux2_1
X_05843_ data_array.rdata0\[4\] net1666 net1147 VGND VGND VPWR VPWR _03356_ sky130_fd_sc_hd__o21a_1
XFILLER_39_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08562_ net707 net4373 net589 VGND VGND VPWR VPWR _00330_ sky130_fd_sc_hd__mux2_1
X_05774_ net9 fsm.tag_out1\[10\] VGND VGND VPWR VPWR _03291_ sky130_fd_sc_hd__nand2_1
XFILLER_35_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07513_ data_array.data1\[5\]\[6\] net1519 net1423 data_array.data1\[6\]\[6\] VGND
+ VGND VPWR VPWR _04748_ sky130_fd_sc_hd__a22o_1
XFILLER_63_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_155_clk clknet_5_28__leaf_clk VGND VGND VPWR VPWR clknet_leaf_155_clk
+ sky130_fd_sc_hd__clkbuf_8
X_08493_ net1711 net626 VGND VGND VPWR VPWR _00293_ sky130_fd_sc_hd__nand2b_1
XFILLER_23_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07444_ data_array.data1\[0\]\[0\] net1366 net1272 data_array.data1\[3\]\[0\] _04684_
+ VGND VGND VPWR VPWR _04685_ sky130_fd_sc_hd__a221o_1
XFILLER_13_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07375_ data_array.data0\[9\]\[58\] net1548 net1452 data_array.data0\[10\]\[58\]
+ VGND VGND VPWR VPWR _04622_ sky130_fd_sc_hd__a22o_1
XFILLER_176_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09114_ net1086 net4326 net566 VGND VGND VPWR VPWR _00868_ sky130_fd_sc_hd__mux2_1
X_06326_ tag_array.tag0\[0\]\[12\] net1402 net1308 tag_array.tag0\[3\]\[12\] _03668_
+ VGND VGND VPWR VPWR _03669_ sky130_fd_sc_hd__a221o_1
X_09045_ net1106 net4091 net410 VGND VGND VPWR VPWR _00799_ sky130_fd_sc_hd__mux2_1
X_06257_ tag_array.tag0\[9\]\[6\] net1564 net1468 tag_array.tag0\[10\]\[6\] VGND VGND
+ VPWR VPWR _03606_ sky130_fd_sc_hd__a22o_1
XFILLER_159_1047 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold430 data_array.data0\[0\]\[30\] VGND VGND VPWR VPWR net2081 sky130_fd_sc_hd__dlygate4sd3_1
X_06188_ tag_array.tag0\[8\]\[0\] net1405 net1311 tag_array.tag0\[11\]\[0\] _03542_
+ VGND VGND VPWR VPWR _03543_ sky130_fd_sc_hd__a221o_1
Xhold441 data_array.data1\[4\]\[5\] VGND VGND VPWR VPWR net2092 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold452 tag_array.tag1\[2\]\[21\] VGND VGND VPWR VPWR net2103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 data_array.data1\[8\]\[3\] VGND VGND VPWR VPWR net2114 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold474 data_array.data0\[4\]\[53\] VGND VGND VPWR VPWR net2125 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold485 data_array.data0\[1\]\[45\] VGND VGND VPWR VPWR net2136 sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 data_array.data1\[10\]\[5\] VGND VGND VPWR VPWR net2147 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_556 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout910 net911 VGND VGND VPWR VPWR net910 sky130_fd_sc_hd__clkbuf_2
XFILLER_132_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_70_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout921 _05514_ VGND VGND VPWR VPWR net921 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout932 _05508_ VGND VGND VPWR VPWR net932 sky130_fd_sc_hd__clkbuf_2
X_09947_ net1042 net3667 net373 VGND VGND VPWR VPWR _01696_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_70_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout943 _05504_ VGND VGND VPWR VPWR net943 sky130_fd_sc_hd__buf_1
XFILLER_89_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout954 _05498_ VGND VGND VPWR VPWR net954 sky130_fd_sc_hd__clkbuf_2
XFILLER_98_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout965 net967 VGND VGND VPWR VPWR net965 sky130_fd_sc_hd__clkbuf_2
XFILLER_58_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout976 net977 VGND VGND VPWR VPWR net976 sky130_fd_sc_hd__clkbuf_2
X_09878_ net956 net4422 net382 VGND VGND VPWR VPWR _01628_ sky130_fd_sc_hd__mux2_1
XFILLER_38_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout987 _05482_ VGND VGND VPWR VPWR net987 sky130_fd_sc_hd__buf_1
XFILLER_135_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout998 net999 VGND VGND VPWR VPWR net998 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_116_Left_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1130 data_array.data1\[2\]\[12\] VGND VGND VPWR VPWR net2781 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1141 data_array.data0\[12\]\[10\] VGND VGND VPWR VPWR net2792 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1152 data_array.data1\[6\]\[5\] VGND VGND VPWR VPWR net2803 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08829_ net1768 net929 net443 VGND VGND VPWR VPWR _00587_ sky130_fd_sc_hd__mux2_1
Xhold1163 tag_array.tag0\[11\]\[4\] VGND VGND VPWR VPWR net2814 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1174 data_array.data1\[12\]\[49\] VGND VGND VPWR VPWR net2825 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1185 data_array.data1\[9\]\[0\] VGND VGND VPWR VPWR net2836 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1196 data_array.data0\[13\]\[34\] VGND VGND VPWR VPWR net2847 sky130_fd_sc_hd__dlygate4sd3_1
X_11840_ clknet_leaf_94_clk _00648_ VGND VGND VPWR VPWR data_array.data0\[7\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_166_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ clknet_leaf_223_clk _00579_ VGND VGND VPWR VPWR data_array.data0\[8\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_68_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_146_clk clknet_5_31__leaf_clk VGND VGND VPWR VPWR clknet_leaf_146_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_26_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13510_ clknet_leaf_83_clk _02139_ VGND VGND VPWR VPWR data_array.data1\[0\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_10722_ net1086 net4420 net490 VGND VGND VPWR VPWR _02467_ sky130_fd_sc_hd__mux2_1
X_14490_ clknet_leaf_101_clk _03113_ VGND VGND VPWR VPWR tag_array.dirty0\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_41_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13441_ clknet_leaf_210_clk _02071_ VGND VGND VPWR VPWR data_array.data1\[8\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10653_ net2008 net1104 net478 VGND VGND VPWR VPWR _02398_ sky130_fd_sc_hd__mux2_1
XFILLER_139_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_125_Left_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13372_ clknet_leaf_109_clk _02002_ VGND VGND VPWR VPWR tag_array.tag0\[2\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_10584_ net871 net2493 net463 VGND VGND VPWR VPWR _02329_ sky130_fd_sc_hd__mux2_1
Xclkload19 clknet_leaf_269_clk VGND VGND VPWR VPWR clkload19/Y sky130_fd_sc_hd__inv_8
XFILLER_6_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12323_ clknet_leaf_202_clk _00055_ VGND VGND VPWR VPWR data_array.rdata0\[5\] sky130_fd_sc_hd__dfxtp_1
X_12254_ clknet_leaf_33_clk _01012_ VGND VGND VPWR VPWR tag_array.tag1\[14\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_182_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11205_ net952 net4589 net649 VGND VGND VPWR VPWR _02948_ sky130_fd_sc_hd__mux2_1
X_12185_ clknet_leaf_108_clk _00993_ VGND VGND VPWR VPWR tag_array.tag0\[14\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11136_ net975 net2263 net543 VGND VGND VPWR VPWR _02879_ sky130_fd_sc_hd__mux2_1
XFILLER_68_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11067_ net2168 net992 net333 VGND VGND VPWR VPWR _02810_ sky130_fd_sc_hd__mux2_1
XFILLER_49_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10018_ net1014 net3399 net563 VGND VGND VPWR VPWR _01767_ sky130_fd_sc_hd__mux2_1
XFILLER_91_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_125_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_125_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11969_ clknet_leaf_47_clk _00777_ VGND VGND VPWR VPWR data_array.data0\[4\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_137_clk clknet_5_31__leaf_clk VGND VGND VPWR VPWR clknet_leaf_137_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13708_ clknet_leaf_69_clk _02337_ VGND VGND VPWR VPWR data_array.data1\[1\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_13639_ clknet_leaf_161_clk _02268_ VGND VGND VPWR VPWR tag_array.dirty0\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_177_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07160_ data_array.data0\[12\]\[38\] net1396 net1302 data_array.data0\[15\]\[38\]
+ _04426_ VGND VGND VPWR VPWR _04427_ sky130_fd_sc_hd__a221o_1
XFILLER_158_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06111_ data_array.rdata0\[26\] net1134 net1113 data_array.rdata1\[26\] VGND VGND
+ VPWR VPWR net281 sky130_fd_sc_hd__a22o_1
X_07091_ data_array.data0\[1\]\[32\] net1526 net1430 data_array.data0\[2\]\[32\] VGND
+ VGND VPWR VPWR _04364_ sky130_fd_sc_hd__a22o_1
X_06042_ fsm.tag_out0\[3\] net1120 _03484_ VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__a21o_1
XFILLER_117_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1031 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_640 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09801_ net1006 net2641 net386 VGND VGND VPWR VPWR _01552_ sky130_fd_sc_hd__mux2_1
XFILLER_113_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07993_ data_array.data1\[5\]\[50\] net1527 net1431 data_array.data1\[6\]\[50\] VGND
+ VGND VPWR VPWR _05184_ sky130_fd_sc_hd__a22o_1
XFILLER_99_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09732_ net760 net4048 net684 VGND VGND VPWR VPWR _01484_ sky130_fd_sc_hd__mux2_1
X_06944_ net1176 _04225_ _04229_ net1224 VGND VGND VPWR VPWR _04231_ sky130_fd_sc_hd__a22o_1
X_09663_ net736 net3045 net612 VGND VGND VPWR VPWR _01415_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06875_ data_array.data0\[5\]\[12\] net1579 net1483 data_array.data0\[6\]\[12\] VGND
+ VGND VPWR VPWR _04168_ sky130_fd_sc_hd__a22o_1
XFILLER_27_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08614_ _05377_ net3006 net518 VGND VGND VPWR VPWR _00373_ sky130_fd_sc_hd__mux2_1
XFILLER_82_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05826_ _03257_ _03260_ _03296_ _03300_ VGND VGND VPWR VPWR _03343_ sky130_fd_sc_hd__or4_1
X_09594_ net973 net3419 net394 VGND VGND VPWR VPWR _01346_ sky130_fd_sc_hd__mux2_1
X_08545_ net774 net3423 net583 VGND VGND VPWR VPWR _00313_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_128_clk clknet_5_30__leaf_clk VGND VGND VPWR VPWR clknet_leaf_128_clk
+ sky130_fd_sc_hd__clkbuf_8
X_05757_ fsm.tag_out1\[13\] net13 VGND VGND VPWR VPWR _03274_ sky130_fd_sc_hd__and2b_1
XFILLER_35_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08476_ net1645 _03146_ VGND VGND VPWR VPWR _05554_ sky130_fd_sc_hd__nor2_1
XFILLER_126_1024 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05688_ fsm.tag_out0\[17\] net17 VGND VGND VPWR VPWR _03205_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_46_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07427_ net1635 _04663_ _04667_ net1209 VGND VGND VPWR VPWR _04670_ sky130_fd_sc_hd__a22o_1
XFILLER_11_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07358_ data_array.data0\[8\]\[56\] net1342 net1248 data_array.data0\[11\]\[56\]
+ _04606_ VGND VGND VPWR VPWR _04607_ sky130_fd_sc_hd__a221o_1
XFILLER_109_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06309_ tag_array.tag0\[12\]\[11\] net1402 net1308 tag_array.tag0\[15\]\[11\] _03652_
+ VGND VGND VPWR VPWR _03653_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_21_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07289_ data_array.data0\[5\]\[50\] net1537 net1441 data_array.data0\[6\]\[50\] VGND
+ VGND VPWR VPWR _04544_ sky130_fd_sc_hd__a22o_1
XFILLER_108_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09028_ net1749 net912 net422 VGND VGND VPWR VPWR _00783_ sky130_fd_sc_hd__mux2_1
XFILLER_151_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_926 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold260 data_array.data0\[2\]\[5\] VGND VGND VPWR VPWR net1911 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold271 tag_array.tag0\[2\]\[21\] VGND VGND VPWR VPWR net1922 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 data_array.data0\[0\]\[19\] VGND VGND VPWR VPWR net1933 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold293 data_array.data0\[1\]\[50\] VGND VGND VPWR VPWR net1944 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_120_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout740 _05391_ VGND VGND VPWR VPWR net740 sky130_fd_sc_hd__clkbuf_2
Xfanout751 net753 VGND VGND VPWR VPWR net751 sky130_fd_sc_hd__clkbuf_2
Xfanout762 net763 VGND VGND VPWR VPWR net762 sky130_fd_sc_hd__clkbuf_2
X_13990_ clknet_leaf_70_clk _02619_ VGND VGND VPWR VPWR data_array.data1\[5\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout773 _05375_ VGND VGND VPWR VPWR net773 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_708 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout784 _05369_ VGND VGND VPWR VPWR net784 sky130_fd_sc_hd__clkbuf_2
Xfanout795 net797 VGND VGND VPWR VPWR net795 sky130_fd_sc_hd__clkbuf_8
X_12941_ clknet_leaf_20_clk _01635_ VGND VGND VPWR VPWR data_array.data0\[13\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_65_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12872_ clknet_leaf_125_clk _01566_ VGND VGND VPWR VPWR data_array.data0\[12\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_142_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11823_ clknet_leaf_268_clk _00631_ VGND VGND VPWR VPWR data_array.data0\[7\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_119_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_119_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_103_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ clknet_leaf_128_clk _00562_ VGND VGND VPWR VPWR data_array.data0\[8\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_83_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10705_ net1821 net898 net479 VGND VGND VPWR VPWR _02450_ sky130_fd_sc_hd__mux2_1
X_14473_ clknet_leaf_249_clk _03096_ VGND VGND VPWR VPWR data_array.data1\[7\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
X_11685_ clknet_leaf_167_clk _00493_ VGND VGND VPWR VPWR tag_array.tag1\[15\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13424_ clknet_leaf_80_clk _02054_ VGND VGND VPWR VPWR data_array.data1\[8\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
X_10636_ net1864 net918 net472 VGND VGND VPWR VPWR _02381_ sky130_fd_sc_hd__mux2_1
Xclkload108 clknet_leaf_34_clk VGND VGND VPWR VPWR clkload108/Y sky130_fd_sc_hd__bufinv_16
Xclkload119 clknet_leaf_75_clk VGND VGND VPWR VPWR clkload119/Y sky130_fd_sc_hd__clkinv_4
X_13355_ clknet_leaf_105_clk _01985_ VGND VGND VPWR VPWR tag_array.tag0\[2\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_10567_ net938 net3540 net460 VGND VGND VPWR VPWR _02312_ sky130_fd_sc_hd__mux2_1
XFILLER_143_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12306_ clknet_leaf_134_clk _01064_ VGND VGND VPWR VPWR tag_array.tag1\[12\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_13286_ clknet_leaf_54_clk _01916_ VGND VGND VPWR VPWR data_array.data0\[11\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
X_10498_ net954 net4146 net345 VGND VGND VPWR VPWR _02243_ sky130_fd_sc_hd__mux2_1
XFILLER_136_990 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_5_14__f_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_5_14__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_5_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12237_ clknet_leaf_145_clk _00166_ VGND VGND VPWR VPWR fsm.tag_out1\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_170_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_3544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12168_ clknet_leaf_160_clk _00976_ VGND VGND VPWR VPWR tag_array.tag0\[14\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_69_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_127_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_3880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11119_ net1040 net2189 net542 VGND VGND VPWR VPWR _02862_ sky130_fd_sc_hd__mux2_1
XFILLER_122_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_127_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12099_ clknet_leaf_28_clk _00907_ VGND VGND VPWR VPWR data_array.data1\[14\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_37_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput6 cpu_addr[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_2
XFILLER_76_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06660_ tag_array.tag1\[13\]\[18\] net1563 net1467 tag_array.tag1\[14\]\[18\] VGND
+ VGND VPWR VPWR _03972_ sky130_fd_sc_hd__a22o_1
XFILLER_92_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06591_ net1629 _03903_ _03907_ net1203 VGND VGND VPWR VPWR _03910_ sky130_fd_sc_hd__a22o_1
XFILLER_51_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08330_ net2102 net1036 net692 VGND VGND VPWR VPWR _00239_ sky130_fd_sc_hd__mux2_1
XFILLER_32_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08261_ fsm.tag_out1\[22\] net816 net808 fsm.tag_out0\[22\] _05408_ VGND VGND VPWR
+ VPWR _05409_ sky130_fd_sc_hd__a221o_2
X_07212_ data_array.data0\[1\]\[43\] net1567 net1471 data_array.data0\[2\]\[43\] VGND
+ VGND VPWR VPWR _04474_ sky130_fd_sc_hd__a22o_1
XFILLER_158_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08192_ _05361_ net815 VGND VGND VPWR VPWR _05362_ sky130_fd_sc_hd__nand2b_1
XFILLER_118_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07143_ _04410_ _04411_ VGND VGND VPWR VPWR _00029_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_41_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07074_ data_array.data0\[0\]\[30\] net1392 net1298 data_array.data0\[3\]\[30\] _04348_
+ VGND VGND VPWR VPWR _04349_ sky130_fd_sc_hd__a221o_1
XFILLER_69_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput310 net310 VGND VGND VPWR VPWR mem_wdata[52] sky130_fd_sc_hd__buf_2
Xoutput321 net321 VGND VGND VPWR VPWR mem_wdata[62] sky130_fd_sc_hd__buf_2
X_06025_ net1162 net23 VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__and2_1
XFILLER_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_929 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07976_ data_array.data1\[0\]\[48\] net1393 net1299 data_array.data1\[3\]\[48\] _05168_
+ VGND VGND VPWR VPWR _05169_ sky130_fd_sc_hd__a221o_1
XFILLER_45_1080 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09715_ net726 net2360 net610 VGND VGND VPWR VPWR _01467_ sky130_fd_sc_hd__mux2_1
X_06927_ data_array.data0\[0\]\[17\] net1336 net1242 data_array.data0\[3\]\[17\] _04214_
+ VGND VGND VPWR VPWR _04215_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_87_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_410 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09646_ net704 net3359 _05571_ VGND VGND VPWR VPWR _01398_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_903 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06858_ data_array.data0\[9\]\[11\] net1568 net1472 data_array.data0\[10\]\[11\]
+ VGND VGND VPWR VPWR _04152_ sky130_fd_sc_hd__a22o_1
XFILLER_27_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_182_Right_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05809_ _03199_ _03321_ _03324_ _03325_ VGND VGND VPWR VPWR _03326_ sky130_fd_sc_hd__or4_1
X_09577_ net1042 net4361 net396 VGND VGND VPWR VPWR _01329_ sky130_fd_sc_hd__mux2_1
XFILLER_55_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06789_ net1630 _04083_ _04087_ net1204 VGND VGND VPWR VPWR _04090_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_65_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08528_ _03507_ _03509_ VGND VGND VPWR VPWR _05590_ sky130_fd_sc_hd__nor2_1
XFILLER_23_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08459_ net1913 net866 net688 VGND VGND VPWR VPWR _00282_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11470_ clknet_leaf_51_clk _00280_ VGND VGND VPWR VPWR data_array.data0\[0\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10421_ net2224 net968 net662 VGND VGND VPWR VPWR _02167_ sky130_fd_sc_hd__mux2_1
XFILLER_109_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13140_ clknet_leaf_32_clk _01834_ VGND VGND VPWR VPWR tag_array.tag1\[8\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_3_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10352_ net794 net3479 net539 VGND VGND VPWR VPWR _02099_ sky130_fd_sc_hd__mux2_1
XFILLER_152_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13071_ clknet_leaf_24_clk _01765_ VGND VGND VPWR VPWR data_array.data1\[13\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_10283_ net3068 net1030 net642 VGND VGND VPWR VPWR _02030_ sky130_fd_sc_hd__mux2_1
XFILLER_183_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12022_ clknet_leaf_264_clk _00830_ VGND VGND VPWR VPWR data_array.data0\[6\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_151_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1502 net1503 VGND VGND VPWR VPWR net1502 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1513 net1516 VGND VGND VPWR VPWR net1513 sky130_fd_sc_hd__clkbuf_4
Xfanout1524 net1543 VGND VGND VPWR VPWR net1524 sky130_fd_sc_hd__buf_2
XFILLER_120_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1535 net1536 VGND VGND VPWR VPWR net1535 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_144_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1546 net1554 VGND VGND VPWR VPWR net1546 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_144_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1557 net1566 VGND VGND VPWR VPWR net1557 sky130_fd_sc_hd__clkbuf_2
Xfanout570 net571 VGND VGND VPWR VPWR net570 sky130_fd_sc_hd__buf_4
XFILLER_93_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1568 net1569 VGND VGND VPWR VPWR net1568 sky130_fd_sc_hd__clkbuf_4
Xfanout581 _05591_ VGND VGND VPWR VPWR net581 sky130_fd_sc_hd__buf_4
XFILLER_76_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1579 net1591 VGND VGND VPWR VPWR net1579 sky130_fd_sc_hd__clkbuf_4
Xfanout592 net594 VGND VGND VPWR VPWR net592 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_161_3452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13973_ clknet_leaf_201_clk _02602_ VGND VGND VPWR VPWR data_array.data1\[5\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_161_3463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12924_ clknet_leaf_31_clk _01618_ VGND VGND VPWR VPWR data_array.data0\[13\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_122_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12855_ clknet_leaf_176_clk _01549_ VGND VGND VPWR VPWR data_array.data0\[12\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11806_ clknet_leaf_16_clk _00614_ VGND VGND VPWR VPWR data_array.data0\[7\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_92_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12786_ clknet_leaf_194_clk _01480_ VGND VGND VPWR VPWR tag_array.tag1\[10\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11737_ clknet_leaf_47_clk _00545_ VGND VGND VPWR VPWR data_array.data0\[8\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_25_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_855 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14456_ clknet_leaf_123_clk _03079_ VGND VGND VPWR VPWR data_array.data1\[7\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_147_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11668_ clknet_leaf_127_clk _00476_ VGND VGND VPWR VPWR tag_array.tag1\[1\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_174_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13407_ clknet_leaf_221_clk _02037_ VGND VGND VPWR VPWR data_array.data1\[8\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_10619_ net2145 net984 net471 VGND VGND VPWR VPWR _02364_ sky130_fd_sc_hd__mux2_1
X_14387_ clknet_leaf_217_clk _03010_ VGND VGND VPWR VPWR data_array.data1\[10\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11599_ clknet_leaf_99_clk _00407_ VGND VGND VPWR VPWR tag_array.tag1\[4\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13338_ clknet_leaf_38_clk _01968_ VGND VGND VPWR VPWR data_array.data0\[10\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_143_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13269_ clknet_leaf_93_clk _01899_ VGND VGND VPWR VPWR data_array.data0\[11\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2408 data_array.data0\[7\]\[6\] VGND VGND VPWR VPWR net4059 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_1012 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_181_3828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2419 data_array.data0\[12\]\[20\] VGND VGND VPWR VPWR net4070 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_181_3839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07830_ data_array.data1\[9\]\[35\] net1525 net1429 data_array.data1\[10\]\[35\]
+ VGND VGND VPWR VPWR _05036_ sky130_fd_sc_hd__a22o_1
Xhold1707 data_array.data1\[11\]\[15\] VGND VGND VPWR VPWR net3358 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1718 data_array.data1\[12\]\[19\] VGND VGND VPWR VPWR net3369 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_99_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1729 data_array.data1\[9\]\[19\] VGND VGND VPWR VPWR net3380 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07761_ data_array.data1\[12\]\[29\] net1387 net1293 data_array.data1\[15\]\[29\]
+ _04972_ VGND VGND VPWR VPWR _04973_ sky130_fd_sc_hd__a221o_1
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09500_ net726 net2446 net626 VGND VGND VPWR VPWR _01253_ sky130_fd_sc_hd__mux2_1
X_06712_ net1196 _04013_ _04017_ net1622 VGND VGND VPWR VPWR _04020_ sky130_fd_sc_hd__a22o_1
XFILLER_53_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07692_ net1217 _04905_ _04909_ net1169 VGND VGND VPWR VPWR _04911_ sky130_fd_sc_hd__a22o_1
XFILLER_25_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09431_ net943 net4579 net587 VGND VGND VPWR VPWR _01184_ sky130_fd_sc_hd__mux2_1
X_06643_ tag_array.tag1\[8\]\[16\] net1417 net1323 tag_array.tag1\[11\]\[16\] _03956_
+ VGND VGND VPWR VPWR _03957_ sky130_fd_sc_hd__a221o_1
XFILLER_92_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09362_ net954 net3951 net405 VGND VGND VPWR VPWR _01115_ sky130_fd_sc_hd__mux2_1
XFILLER_24_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06574_ tag_array.tag1\[1\]\[10\] net1595 net1499 tag_array.tag1\[2\]\[10\] VGND
+ VGND VPWR VPWR _03894_ sky130_fd_sc_hd__a22o_1
XFILLER_33_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08313_ net103 net38 net1644 VGND VGND VPWR VPWR _05445_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09293_ net706 net2644 net563 VGND VGND VPWR VPWR _01047_ sky130_fd_sc_hd__mux2_1
XANTENNA_11 _00173_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_22 _03513_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08244_ net729 net4479 net804 VGND VGND VPWR VPWR _00212_ sky130_fd_sc_hd__mux2_1
XANTENNA_33 net340 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_44 net556 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_55 net1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_66 net1627 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_77 net369 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08175_ net1201 _05343_ _05347_ net1626 VGND VGND VPWR VPWR _05350_ sky130_fd_sc_hd__a22o_1
XANTENNA_88 net1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07126_ data_array.data0\[9\]\[35\] net1537 net1441 data_array.data0\[10\]\[35\]
+ VGND VGND VPWR VPWR _04396_ sky130_fd_sc_hd__a22o_1
XFILLER_174_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07057_ data_array.data0\[12\]\[29\] net1380 net1286 data_array.data0\[15\]\[29\]
+ _04332_ VGND VGND VPWR VPWR _04333_ sky130_fd_sc_hd__a221o_1
XFILLER_115_960 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06008_ data_array.rdata0\[59\] net1658 net1148 VGND VGND VPWR VPWR _03466_ sky130_fd_sc_hd__o21a_1
Xoutput173 net173 VGND VGND VPWR VPWR cpu_rdata[17] sky130_fd_sc_hd__buf_2
XFILLER_115_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput184 net184 VGND VGND VPWR VPWR cpu_rdata[27] sky130_fd_sc_hd__clkbuf_4
Xoutput195 net195 VGND VGND VPWR VPWR cpu_rdata[37] sky130_fd_sc_hd__clkbuf_4
Xhold2920 data_array.data1\[10\]\[48\] VGND VGND VPWR VPWR net4571 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2931 data_array.data0\[11\]\[26\] VGND VGND VPWR VPWR net4582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2942 data_array.data1\[15\]\[9\] VGND VGND VPWR VPWR net4593 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2953 tag_array.tag0\[6\]\[7\] VGND VGND VPWR VPWR net4604 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2964 data_array.data0\[7\]\[1\] VGND VGND VPWR VPWR net4615 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2975 net327 VGND VGND VPWR VPWR net4626 sky130_fd_sc_hd__dlygate4sd3_1
X_07959_ data_array.data1\[8\]\[47\] net1397 net1303 data_array.data1\[11\]\[47\]
+ _05152_ VGND VGND VPWR VPWR _05153_ sky130_fd_sc_hd__a221o_1
XFILLER_75_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10970_ net862 net3265 net535 VGND VGND VPWR VPWR _02715_ sky130_fd_sc_hd__mux2_1
XFILLER_55_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09629_ net771 net3260 net617 VGND VGND VPWR VPWR _01381_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_100_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12640_ clknet_leaf_22_clk _01334_ VGND VGND VPWR VPWR data_array.data0\[15\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_80_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12571_ clknet_leaf_171_clk _01265_ VGND VGND VPWR VPWR tag_array.tag0\[10\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_50_clk clknet_5_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_50_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_184_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14310_ clknet_leaf_67_clk _02939_ VGND VGND VPWR VPWR data_array.data1\[11\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11522_ clknet_leaf_102_clk _00330_ VGND VGND VPWR VPWR tag_array.tag1\[9\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_178_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14241_ clknet_leaf_263_clk _02870_ VGND VGND VPWR VPWR data_array.data1\[12\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11453_ clknet_leaf_93_clk _00263_ VGND VGND VPWR VPWR data_array.data0\[0\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10404_ net2433 net1038 net667 VGND VGND VPWR VPWR _02150_ sky130_fd_sc_hd__mux2_1
X_14172_ clknet_leaf_125_clk _02801_ VGND VGND VPWR VPWR data_array.data0\[2\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_11384_ net164 VGND VGND VPWR VPWR _00194_ sky130_fd_sc_hd__inv_2
XFILLER_178_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13123_ clknet_leaf_105_clk _01817_ VGND VGND VPWR VPWR tag_array.tag0\[3\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_10335_ net758 net3396 net592 VGND VGND VPWR VPWR _02082_ sky130_fd_sc_hd__mux2_1
XFILLER_11_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13054_ clknet_leaf_197_clk _01748_ VGND VGND VPWR VPWR data_array.data1\[13\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_112_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_163_3503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10266_ net2114 net1099 net635 VGND VGND VPWR VPWR _02013_ sky130_fd_sc_hd__mux2_1
XFILLER_97_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12005_ clknet_leaf_63_clk _00813_ VGND VGND VPWR VPWR data_array.data0\[6\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout1310 net1312 VGND VGND VPWR VPWR net1310 sky130_fd_sc_hd__clkbuf_4
Xfanout1321 net1322 VGND VGND VPWR VPWR net1321 sky130_fd_sc_hd__clkbuf_4
Xfanout1332 net1334 VGND VGND VPWR VPWR net1332 sky130_fd_sc_hd__clkbuf_4
X_10197_ net1019 net3818 net356 VGND VGND VPWR VPWR _01944_ sky130_fd_sc_hd__mux2_1
XFILLER_66_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1343 net1345 VGND VGND VPWR VPWR net1343 sky130_fd_sc_hd__clkbuf_4
XFILLER_121_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1354 net1355 VGND VGND VPWR VPWR net1354 sky130_fd_sc_hd__clkbuf_4
Xfanout1365 net1367 VGND VGND VPWR VPWR net1365 sky130_fd_sc_hd__clkbuf_4
Xfanout1376 _03513_ VGND VGND VPWR VPWR net1376 sky130_fd_sc_hd__buf_4
XFILLER_78_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1387 net1388 VGND VGND VPWR VPWR net1387 sky130_fd_sc_hd__clkbuf_4
Xfanout1398 net1399 VGND VGND VPWR VPWR net1398 sky130_fd_sc_hd__clkbuf_4
XFILLER_4_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13956_ clknet_leaf_120_clk _02585_ VGND VGND VPWR VPWR data_array.data1\[4\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12907_ clknet_leaf_45_clk _01601_ VGND VGND VPWR VPWR data_array.data0\[13\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_13887_ clknet_leaf_17_clk _02516_ VGND VGND VPWR VPWR data_array.data1\[3\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
X_12838_ clknet_leaf_0_clk _01532_ VGND VGND VPWR VPWR data_array.data0\[12\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12769_ clknet_leaf_155_clk _01463_ VGND VGND VPWR VPWR tag_array.tag0\[6\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_41_clk clknet_5_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_41_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_175_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06290_ tag_array.tag0\[9\]\[9\] net1598 net1502 tag_array.tag0\[10\]\[9\] VGND VGND
+ VPWR VPWR _03636_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_174_3698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput20 cpu_addr[27] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_2
X_14439_ clknet_leaf_203_clk _03062_ VGND VGND VPWR VPWR data_array.data1\[7\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput31 cpu_addr[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_135_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput42 cpu_wdata[17] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_1
Xinput53 cpu_wdata[27] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_1
XFILLER_116_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput64 cpu_wdata[37] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput75 cpu_wdata[47] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_1
Xhold804 data_array.data1\[2\]\[47\] VGND VGND VPWR VPWR net2455 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_156_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput86 cpu_wdata[57] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_1
Xhold815 tag_array.tag0\[2\]\[19\] VGND VGND VPWR VPWR net2466 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold826 data_array.data0\[3\]\[29\] VGND VGND VPWR VPWR net2477 sky130_fd_sc_hd__dlygate4sd3_1
Xinput97 cpu_wdata[9] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_1
Xhold837 data_array.data0\[9\]\[49\] VGND VGND VPWR VPWR net2488 sky130_fd_sc_hd__dlygate4sd3_1
Xhold848 data_array.data1\[13\]\[34\] VGND VGND VPWR VPWR net2499 sky130_fd_sc_hd__dlygate4sd3_1
X_09980_ net909 net3814 net371 VGND VGND VPWR VPWR _01729_ sky130_fd_sc_hd__mux2_1
Xhold859 tag_array.tag1\[6\]\[1\] VGND VGND VPWR VPWR net2510 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08931_ net1042 net4021 net428 VGND VGND VPWR VPWR _00687_ sky130_fd_sc_hd__mux2_1
XFILLER_103_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2205 data_array.data0\[13\]\[51\] VGND VGND VPWR VPWR net3856 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2216 data_array.data0\[6\]\[59\] VGND VGND VPWR VPWR net3867 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_36_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08862_ net1058 net3976 net436 VGND VGND VPWR VPWR _00619_ sky130_fd_sc_hd__mux2_1
Xhold2227 tag_array.tag0\[11\]\[9\] VGND VGND VPWR VPWR net3878 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_36_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2238 data_array.data1\[13\]\[22\] VGND VGND VPWR VPWR net3889 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2249 data_array.data1\[3\]\[41\] VGND VGND VPWR VPWR net3900 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1504 tag_array.tag0\[11\]\[18\] VGND VGND VPWR VPWR net3155 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1515 data_array.data0\[3\]\[31\] VGND VGND VPWR VPWR net3166 sky130_fd_sc_hd__dlygate4sd3_1
X_07813_ net1228 _05015_ _05019_ net1180 VGND VGND VPWR VPWR _05021_ sky130_fd_sc_hd__a22o_1
Xhold1526 tag_array.tag0\[13\]\[14\] VGND VGND VPWR VPWR net3177 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1537 data_array.data1\[7\]\[21\] VGND VGND VPWR VPWR net3188 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08793_ net1772 net1073 net447 VGND VGND VPWR VPWR _00551_ sky130_fd_sc_hd__mux2_1
Xhold1548 data_array.data1\[11\]\[37\] VGND VGND VPWR VPWR net3199 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1559 data_array.data0\[15\]\[27\] VGND VGND VPWR VPWR net3210 sky130_fd_sc_hd__dlygate4sd3_1
X_07744_ data_array.data1\[5\]\[27\] net1547 net1451 data_array.data1\[6\]\[27\] VGND
+ VGND VPWR VPWR _04958_ sky130_fd_sc_hd__a22o_1
XFILLER_25_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07675_ data_array.data1\[0\]\[21\] net1365 net1271 data_array.data1\[3\]\[21\] _04894_
+ VGND VGND VPWR VPWR _04895_ sky130_fd_sc_hd__a221o_1
XFILLER_65_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09414_ net1008 net4154 net578 VGND VGND VPWR VPWR _01167_ sky130_fd_sc_hd__mux2_1
X_06626_ _03940_ _03941_ VGND VGND VPWR VPWR _00161_ sky130_fd_sc_hd__or2_2
X_09345_ net1020 net4175 net403 VGND VGND VPWR VPWR _01098_ sky130_fd_sc_hd__mux2_1
XFILLER_80_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06557_ tag_array.tag1\[0\]\[8\] net1417 net1323 tag_array.tag1\[3\]\[8\] _03878_
+ VGND VGND VPWR VPWR _03879_ sky130_fd_sc_hd__a221o_1
XFILLER_139_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_32_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_21_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09276_ net774 net3538 net558 VGND VGND VPWR VPWR _01030_ sky130_fd_sc_hd__mux2_1
X_06488_ tag_array.tag1\[13\]\[2\] net1541 net1445 tag_array.tag1\[14\]\[2\] VGND
+ VGND VPWR VPWR _03816_ sky130_fd_sc_hd__a22o_1
XFILLER_138_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08227_ _03139_ _03147_ VGND VGND VPWR VPWR _05386_ sky130_fd_sc_hd__nor2_1
XFILLER_138_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08158_ tag_array.dirty0\[1\] net1594 net1498 tag_array.dirty0\[2\] VGND VGND VPWR
+ VPWR _05334_ sky130_fd_sc_hd__a22o_1
XFILLER_146_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07109_ net1227 _04375_ _04379_ net1179 VGND VGND VPWR VPWR _04381_ sky130_fd_sc_hd__a22o_1
X_08089_ _05270_ _05271_ VGND VGND VPWR VPWR _00117_ sky130_fd_sc_hd__or2_1
XFILLER_134_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10120_ net1065 net4441 net366 VGND VGND VPWR VPWR _01868_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_99_clk clknet_5_24__leaf_clk VGND VGND VPWR VPWR clknet_leaf_99_clk sky130_fd_sc_hd__clkbuf_8
X_10051_ net882 net3652 net555 VGND VGND VPWR VPWR _01800_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_73_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2750 data_array.data1\[14\]\[47\] VGND VGND VPWR VPWR net4401 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2761 data_array.data1\[6\]\[43\] VGND VGND VPWR VPWR net4412 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2772 tag_array.tag1\[9\]\[12\] VGND VGND VPWR VPWR net4423 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_169_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2783 data_array.data1\[7\]\[9\] VGND VGND VPWR VPWR net4434 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_169_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2794 data_array.data0\[13\]\[24\] VGND VGND VPWR VPWR net4445 sky130_fd_sc_hd__dlygate4sd3_1
X_13810_ clknet_leaf_88_clk _02439_ VGND VGND VPWR VPWR data_array.data1\[2\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13741_ clknet_leaf_214_clk _02370_ VGND VGND VPWR VPWR data_array.data1\[1\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_27_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10953_ net930 net4477 net530 VGND VGND VPWR VPWR _02698_ sky130_fd_sc_hd__mux2_1
XFILLER_16_446 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13672_ clknet_leaf_258_clk _02301_ VGND VGND VPWR VPWR data_array.data1\[15\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
X_10884_ net950 net4340 net523 VGND VGND VPWR VPWR _02629_ sky130_fd_sc_hd__mux2_1
XFILLER_73_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_139_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12623_ clknet_leaf_203_clk _01317_ VGND VGND VPWR VPWR data_array.data0\[15\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_1052 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_23_clk clknet_5_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_156_3362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12554_ clknet_leaf_161_clk _01248_ VGND VGND VPWR VPWR tag_array.tag0\[11\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11505_ clknet_leaf_196_clk _00313_ VGND VGND VPWR VPWR tag_array.tag1\[9\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_117_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12485_ clknet_leaf_213_clk _01179_ VGND VGND VPWR VPWR data_array.data1\[9\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_172_616 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14224_ clknet_leaf_19_clk _02853_ VGND VGND VPWR VPWR data_array.data1\[12\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_11436_ clknet_leaf_263_clk _00246_ VGND VGND VPWR VPWR data_array.data0\[0\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_153_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14155_ clknet_leaf_48_clk _02784_ VGND VGND VPWR VPWR data_array.data0\[2\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_11367_ net1646 net4312 net610 VGND VGND VPWR VPWR _03110_ sky130_fd_sc_hd__mux2_1
X_13106_ clknet_leaf_239_clk _01800_ VGND VGND VPWR VPWR data_array.data1\[13\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_130_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10318_ net1994 net890 net635 VGND VGND VPWR VPWR _02065_ sky130_fd_sc_hd__mux2_1
XFILLER_112_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14086_ clknet_leaf_120_clk _02715_ VGND VGND VPWR VPWR data_array.data1\[6\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11298_ net1100 net2216 net797 VGND VGND VPWR VPWR _03041_ sky130_fd_sc_hd__mux2_1
XFILLER_65_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13037_ clknet_leaf_223_clk _01731_ VGND VGND VPWR VPWR data_array.data0\[3\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10249_ net748 net3336 net596 VGND VGND VPWR VPWR _01996_ sky130_fd_sc_hd__mux2_1
Xfanout1140 net1141 VGND VGND VPWR VPWR net1140 sky130_fd_sc_hd__buf_4
XFILLER_26_1067 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1151 net1154 VGND VGND VPWR VPWR net1151 sky130_fd_sc_hd__buf_4
Xfanout1162 net262 VGND VGND VPWR VPWR net1162 sky130_fd_sc_hd__clkbuf_2
XFILLER_66_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1173 net1174 VGND VGND VPWR VPWR net1173 sky130_fd_sc_hd__buf_4
Xfanout1184 net1186 VGND VGND VPWR VPWR net1184 sky130_fd_sc_hd__clkbuf_4
Xfanout1195 net1198 VGND VGND VPWR VPWR net1195 sky130_fd_sc_hd__buf_4
XFILLER_82_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05790_ _03283_ _03304_ _03305_ _03306_ VGND VGND VPWR VPWR _03307_ sky130_fd_sc_hd__or4_1
XFILLER_81_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13939_ clknet_leaf_44_clk _02568_ VGND VGND VPWR VPWR data_array.data1\[4\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_755 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_176_3738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07460_ net1188 _04693_ _04697_ net1614 VGND VGND VPWR VPWR _04700_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_176_3749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06411_ tag_array.tag0\[9\]\[20\] net1559 net1463 tag_array.tag0\[10\]\[20\] VGND
+ VGND VPWR VPWR _03746_ sky130_fd_sc_hd__a22o_1
X_07391_ data_array.data0\[12\]\[59\] net1379 net1285 data_array.data0\[15\]\[59\]
+ _04636_ VGND VGND VPWR VPWR _04637_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_14_clk clknet_5_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_8
X_09130_ net1021 net3025 net568 VGND VGND VPWR VPWR _00884_ sky130_fd_sc_hd__mux2_1
X_06342_ tag_array.tag0\[8\]\[14\] net1369 net1275 tag_array.tag0\[11\]\[14\] _03682_
+ VGND VGND VPWR VPWR _03683_ sky130_fd_sc_hd__a221o_1
X_09061_ net1042 net3332 net412 VGND VGND VPWR VPWR _00815_ sky130_fd_sc_hd__mux2_1
X_06273_ net1232 _03615_ _03619_ net1184 VGND VGND VPWR VPWR _03621_ sky130_fd_sc_hd__a22o_1
XFILLER_175_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08012_ _05200_ _05201_ VGND VGND VPWR VPWR _00110_ sky130_fd_sc_hd__or2_1
Xhold601 data_array.data1\[0\]\[30\] VGND VGND VPWR VPWR net2252 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold612 data_array.data1\[12\]\[34\] VGND VGND VPWR VPWR net2263 sky130_fd_sc_hd__dlygate4sd3_1
Xhold623 data_array.data0\[4\]\[27\] VGND VGND VPWR VPWR net2274 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold634 tag_array.tag1\[10\]\[18\] VGND VGND VPWR VPWR net2285 sky130_fd_sc_hd__dlygate4sd3_1
Xhold645 tag_array.tag1\[2\]\[23\] VGND VGND VPWR VPWR net2296 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold656 data_array.data0\[14\]\[37\] VGND VGND VPWR VPWR net2307 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold667 data_array.data0\[8\]\[51\] VGND VGND VPWR VPWR net2318 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold678 tag_array.tag1\[7\]\[4\] VGND VGND VPWR VPWR net2329 sky130_fd_sc_hd__dlygate4sd3_1
X_09963_ net976 net4244 net375 VGND VGND VPWR VPWR _01712_ sky130_fd_sc_hd__mux2_1
Xhold689 data_array.data1\[5\]\[17\] VGND VGND VPWR VPWR net2340 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2002 data_array.data1\[10\]\[37\] VGND VGND VPWR VPWR net3653 sky130_fd_sc_hd__dlygate4sd3_1
X_08914_ net1108 net3353 net429 VGND VGND VPWR VPWR _00670_ sky130_fd_sc_hd__mux2_1
Xhold2013 tag_array.tag0\[7\]\[18\] VGND VGND VPWR VPWR net3664 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09894_ net894 net4107 net380 VGND VGND VPWR VPWR _01644_ sky130_fd_sc_hd__mux2_1
Xhold2024 data_array.data0\[5\]\[23\] VGND VGND VPWR VPWR net3675 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2035 tag_array.tag0\[5\]\[11\] VGND VGND VPWR VPWR net3686 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2046 data_array.data1\[10\]\[11\] VGND VGND VPWR VPWR net3697 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1301 data_array.data0\[5\]\[48\] VGND VGND VPWR VPWR net2952 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2057 data_array.data1\[6\]\[63\] VGND VGND VPWR VPWR net3708 sky130_fd_sc_hd__dlygate4sd3_1
X_08845_ net2187 net867 net445 VGND VGND VPWR VPWR _00603_ sky130_fd_sc_hd__mux2_1
Xhold1312 tag_array.tag0\[3\]\[18\] VGND VGND VPWR VPWR net2963 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2068 data_array.data1\[5\]\[62\] VGND VGND VPWR VPWR net3719 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_40_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_51_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1323 tag_array.tag0\[14\]\[3\] VGND VGND VPWR VPWR net2974 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1334 data_array.data1\[5\]\[54\] VGND VGND VPWR VPWR net2985 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2079 data_array.data0\[7\]\[9\] VGND VGND VPWR VPWR net3730 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1345 tag_array.tag0\[13\]\[6\] VGND VGND VPWR VPWR net2996 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1356 data_array.data0\[3\]\[25\] VGND VGND VPWR VPWR net3007 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1367 data_array.data0\[4\]\[4\] VGND VGND VPWR VPWR net3018 sky130_fd_sc_hd__dlygate4sd3_1
X_08776_ net719 net3450 net450 VGND VGND VPWR VPWR _00535_ sky130_fd_sc_hd__mux2_1
X_05988_ data_array.rdata1\[52\] net830 net839 VGND VGND VPWR VPWR _03453_ sky130_fd_sc_hd__a21o_1
Xhold1378 data_array.data0\[10\]\[39\] VGND VGND VPWR VPWR net3029 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1389 tag_array.tag1\[15\]\[6\] VGND VGND VPWR VPWR net3040 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07727_ data_array.data1\[9\]\[26\] net1525 net1429 data_array.data1\[10\]\[26\]
+ VGND VGND VPWR VPWR _04942_ sky130_fd_sc_hd__a22o_1
XFILLER_27_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07658_ net1206 _04873_ _04877_ net1632 VGND VGND VPWR VPWR _04880_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06609_ tag_array.tag1\[9\]\[13\] net1611 net1515 tag_array.tag1\[10\]\[13\] VGND
+ VGND VPWR VPWR _03926_ sky130_fd_sc_hd__a22o_1
XFILLER_43_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07589_ data_array.data1\[8\]\[13\] net1364 net1270 data_array.data1\[11\]\[13\]
+ _04816_ VGND VGND VPWR VPWR _04817_ sky130_fd_sc_hd__a221o_1
XFILLER_13_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_8_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_8_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_139_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09328_ net1088 net2386 net404 VGND VGND VPWR VPWR _01081_ sky130_fd_sc_hd__mux2_1
XFILLER_159_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09259_ net742 net3057 net571 VGND VGND VPWR VPWR _01013_ sky130_fd_sc_hd__mux2_1
XFILLER_182_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12270_ clknet_leaf_31_clk _01028_ VGND VGND VPWR VPWR tag_array.tag1\[13\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_138_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11221_ net891 net4014 net650 VGND VGND VPWR VPWR _02964_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_112_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11152_ net911 net3917 net541 VGND VGND VPWR VPWR _02895_ sky130_fd_sc_hd__mux2_1
XFILLER_49_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10103_ net4215 net711 net636 VGND VGND VPWR VPWR _01852_ sky130_fd_sc_hd__mux2_1
XFILLER_0_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11083_ net2904 net928 net329 VGND VGND VPWR VPWR _02826_ sky130_fd_sc_hd__mux2_1
X_10034_ net951 net3993 net564 VGND VGND VPWR VPWR _01783_ sky130_fd_sc_hd__mux2_1
Xhold2580 data_array.data1\[10\]\[43\] VGND VGND VPWR VPWR net4231 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2591 data_array.data1\[12\]\[46\] VGND VGND VPWR VPWR net4242 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_124_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1890 data_array.data1\[10\]\[19\] VGND VGND VPWR VPWR net3541 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11985_ clknet_leaf_52_clk _00793_ VGND VGND VPWR VPWR data_array.data0\[4\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_158_3402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13724_ clknet_leaf_122_clk _02353_ VGND VGND VPWR VPWR data_array.data1\[1\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_10936_ net996 net4039 net530 VGND VGND VPWR VPWR _02681_ sky130_fd_sc_hd__mux2_1
XFILLER_140_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13655_ clknet_leaf_70_clk _02284_ VGND VGND VPWR VPWR data_array.data1\[15\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_10867_ net1017 net3077 net516 VGND VGND VPWR VPWR _02612_ sky130_fd_sc_hd__mux2_1
XFILLER_32_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12606_ clknet_leaf_138_clk _01300_ VGND VGND VPWR VPWR tag_array.tag0\[0\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13586_ clknet_leaf_45_clk _02215_ VGND VGND VPWR VPWR data_array.data0\[9\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_169_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10798_ net2033 net1038 net503 VGND VGND VPWR VPWR _02543_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_171_3646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12537_ clknet_leaf_102_clk _01231_ VGND VGND VPWR VPWR tag_array.tag1\[11\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_30_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_132_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12468_ clknet_leaf_122_clk _01162_ VGND VGND VPWR VPWR data_array.data1\[9\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14207_ clknet_leaf_14_clk _02836_ VGND VGND VPWR VPWR data_array.data0\[2\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
X_11419_ clknet_leaf_16_clk _00229_ VGND VGND VPWR VPWR data_array.data0\[0\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_12399_ clknet_leaf_246_clk _01093_ VGND VGND VPWR VPWR data_array.data0\[14\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_153_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14138_ clknet_leaf_241_clk _02767_ VGND VGND VPWR VPWR data_array.data0\[1\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06960_ data_array.data0\[4\]\[20\] net1413 net1319 data_array.data0\[7\]\[20\] _04244_
+ VGND VGND VPWR VPWR _04245_ sky130_fd_sc_hd__a221o_1
X_14069_ clknet_leaf_26_clk _02698_ VGND VGND VPWR VPWR data_array.data1\[6\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_579 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_3_clk clknet_5_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_33_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05911_ net117 net1150 _03400_ _03401_ VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__a22o_1
XFILLER_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06891_ data_array.data0\[9\]\[14\] net1569 net1473 data_array.data0\[10\]\[14\]
+ VGND VGND VPWR VPWR _04182_ sky130_fd_sc_hd__a22o_1
X_08630_ net703 net2389 net516 VGND VGND VPWR VPWR _00389_ sky130_fd_sc_hd__mux2_1
XFILLER_95_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05842_ net132 net1156 _03355_ _03354_ VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__a22o_1
XFILLER_54_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08561_ net710 net4398 net580 VGND VGND VPWR VPWR _00329_ sky130_fd_sc_hd__mux2_1
XFILLER_82_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05773_ _03247_ _03248_ _03289_ VGND VGND VPWR VPWR _03290_ sky130_fd_sc_hd__or3_1
X_07512_ data_array.data1\[12\]\[6\] net1329 net1235 data_array.data1\[15\]\[6\] _04746_
+ VGND VGND VPWR VPWR _04747_ sky130_fd_sc_hd__a221o_1
XFILLER_81_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08492_ net825 net815 _05550_ net855 VGND VGND VPWR VPWR _05565_ sky130_fd_sc_hd__or4_4
XFILLER_120_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_736 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07443_ data_array.data1\[1\]\[0\] net1556 net1460 data_array.data1\[2\]\[0\] VGND
+ VGND VPWR VPWR _04684_ sky130_fd_sc_hd__a22o_1
XFILLER_90_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07374_ _04620_ _04621_ VGND VGND VPWR VPWR _00052_ sky130_fd_sc_hd__or2_1
XFILLER_148_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09113_ net1091 net4209 net570 VGND VGND VPWR VPWR _00867_ sky130_fd_sc_hd__mux2_1
X_06325_ tag_array.tag0\[1\]\[12\] net1593 net1497 tag_array.tag0\[2\]\[12\] VGND
+ VGND VPWR VPWR _03668_ sky130_fd_sc_hd__a22o_1
XFILLER_129_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_616 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09044_ net1108 net3411 net413 VGND VGND VPWR VPWR _00798_ sky130_fd_sc_hd__mux2_1
X_06256_ tag_array.tag0\[4\]\[6\] net1373 net1279 tag_array.tag0\[7\]\[6\] _03604_
+ VGND VGND VPWR VPWR _03605_ sky130_fd_sc_hd__a221o_1
XFILLER_117_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold420 data_array.data1\[2\]\[5\] VGND VGND VPWR VPWR net2071 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold431 data_array.data0\[1\]\[26\] VGND VGND VPWR VPWR net2082 sky130_fd_sc_hd__dlygate4sd3_1
X_06187_ tag_array.tag0\[9\]\[0\] net1596 net1500 tag_array.tag0\[10\]\[0\] VGND VGND
+ VPWR VPWR _03542_ sky130_fd_sc_hd__a22o_1
Xhold442 data_array.data1\[2\]\[54\] VGND VGND VPWR VPWR net2093 sky130_fd_sc_hd__dlygate4sd3_1
Xhold453 data_array.data1\[4\]\[62\] VGND VGND VPWR VPWR net2104 sky130_fd_sc_hd__dlygate4sd3_1
Xhold464 tag_array.tag1\[10\]\[22\] VGND VGND VPWR VPWR net2115 sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 data_array.data0\[3\]\[15\] VGND VGND VPWR VPWR net2126 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold486 data_array.data0\[1\]\[9\] VGND VGND VPWR VPWR net2137 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout900 _05524_ VGND VGND VPWR VPWR net900 sky130_fd_sc_hd__clkbuf_2
XFILLER_132_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout911 _05520_ VGND VGND VPWR VPWR net911 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold497 data_array.data1\[4\]\[24\] VGND VGND VPWR VPWR net2148 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout922 net923 VGND VGND VPWR VPWR net922 sky130_fd_sc_hd__clkbuf_2
XFILLER_77_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09946_ net1046 net3781 net373 VGND VGND VPWR VPWR _01695_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_70_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout933 _05508_ VGND VGND VPWR VPWR net933 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_70_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout944 net947 VGND VGND VPWR VPWR net944 sky130_fd_sc_hd__clkbuf_2
Xfanout955 _05498_ VGND VGND VPWR VPWR net955 sky130_fd_sc_hd__buf_1
XFILLER_86_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout966 net967 VGND VGND VPWR VPWR net966 sky130_fd_sc_hd__clkbuf_2
Xfanout977 net979 VGND VGND VPWR VPWR net977 sky130_fd_sc_hd__clkbuf_2
X_09877_ net961 net2650 net380 VGND VGND VPWR VPWR _01627_ sky130_fd_sc_hd__mux2_1
XFILLER_57_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1120 tag_array.tag0\[8\]\[1\] VGND VGND VPWR VPWR net2771 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout988 net989 VGND VGND VPWR VPWR net988 sky130_fd_sc_hd__clkbuf_2
Xfanout999 _05476_ VGND VGND VPWR VPWR net999 sky130_fd_sc_hd__buf_1
XFILLER_100_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1131 data_array.data1\[13\]\[31\] VGND VGND VPWR VPWR net2782 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1142 tag_array.tag1\[3\]\[6\] VGND VGND VPWR VPWR net2793 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08828_ net2087 net933 net448 VGND VGND VPWR VPWR _00586_ sky130_fd_sc_hd__mux2_1
Xhold1153 data_array.data0\[11\]\[63\] VGND VGND VPWR VPWR net2804 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_161_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1164 data_array.data1\[9\]\[9\] VGND VGND VPWR VPWR net2815 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1175 data_array.data1\[0\]\[51\] VGND VGND VPWR VPWR net2826 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_79_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1186 data_array.data0\[0\]\[20\] VGND VGND VPWR VPWR net2837 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08759_ net790 net3274 net450 VGND VGND VPWR VPWR _00518_ sky130_fd_sc_hd__mux2_1
Xhold1197 tag_array.tag0\[13\]\[12\] VGND VGND VPWR VPWR net2848 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_16_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ clknet_leaf_114_clk _00578_ VGND VGND VPWR VPWR data_array.data0\[8\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_41_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ net1090 net3597 net493 VGND VGND VPWR VPWR _02466_ sky130_fd_sc_hd__mux2_1
X_13440_ clknet_leaf_120_clk _02070_ VGND VGND VPWR VPWR data_array.data1\[8\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_153_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10652_ net2227 net1110 net482 VGND VGND VPWR VPWR _02397_ sky130_fd_sc_hd__mux2_1
XFILLER_41_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13371_ clknet_leaf_157_clk _02001_ VGND VGND VPWR VPWR tag_array.tag0\[2\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_155_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10583_ net875 net3322 net460 VGND VGND VPWR VPWR _02328_ sky130_fd_sc_hd__mux2_1
XFILLER_103_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12322_ clknet_leaf_76_clk _00044_ VGND VGND VPWR VPWR data_array.rdata0\[4\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_88_Right_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12253_ clknet_leaf_105_clk _01011_ VGND VGND VPWR VPWR tag_array.tag1\[14\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_108_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11204_ net959 net4572 net656 VGND VGND VPWR VPWR _02947_ sky130_fd_sc_hd__mux2_1
XFILLER_79_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12184_ clknet_leaf_157_clk _00992_ VGND VGND VPWR VPWR tag_array.tag0\[14\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11135_ net978 net3086 net549 VGND VGND VPWR VPWR _02878_ sky130_fd_sc_hd__mux2_1
XFILLER_123_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11066_ net1970 net996 net329 VGND VGND VPWR VPWR _02809_ sky130_fd_sc_hd__mux2_1
XFILLER_77_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10017_ net1016 net3561 net558 VGND VGND VPWR VPWR _01766_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_97_Right_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_125_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11968_ clknet_leaf_96_clk _00776_ VGND VGND VPWR VPWR data_array.data0\[4\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_45_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13707_ clknet_leaf_36_clk _02336_ VGND VGND VPWR VPWR data_array.data1\[1\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_10919_ net1067 net3810 net534 VGND VGND VPWR VPWR _02664_ sky130_fd_sc_hd__mux2_1
X_11899_ clknet_leaf_216_clk _00707_ VGND VGND VPWR VPWR data_array.data0\[5\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_71_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13638_ clknet_leaf_224_clk _02267_ VGND VGND VPWR VPWR data_array.data0\[9\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
X_13569_ clknet_leaf_29_clk _02198_ VGND VGND VPWR VPWR tag_array.dirty1\[5\] sky130_fd_sc_hd__dfxtp_1
X_06110_ data_array.rdata0\[25\] net1134 net1112 data_array.rdata1\[25\] VGND VGND
+ VPWR VPWR net280 sky130_fd_sc_hd__a22o_1
X_07090_ data_array.data0\[12\]\[32\] net1333 net1239 data_array.data0\[15\]\[32\]
+ _04362_ VGND VGND VPWR VPWR _04363_ sky130_fd_sc_hd__a221o_1
XFILLER_172_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06041_ net1158 net2 fsm.tag_out1\[3\] net1131 VGND VGND VPWR VPWR _03484_ sky130_fd_sc_hd__a22o_1
XFILLER_114_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_1043 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09800_ net1010 net2986 net386 VGND VGND VPWR VPWR _01551_ sky130_fd_sc_hd__mux2_1
X_07992_ data_array.data1\[8\]\[50\] net1346 net1252 data_array.data1\[11\]\[50\]
+ _05182_ VGND VGND VPWR VPWR _05183_ sky130_fd_sc_hd__a221o_1
X_09731_ net765 net2501 net683 VGND VGND VPWR VPWR _01483_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_163_Right_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06943_ net1618 _04223_ _04227_ net1192 VGND VGND VPWR VPWR _04230_ sky130_fd_sc_hd__a22o_1
XFILLER_86_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09662_ net738 net2374 net613 VGND VGND VPWR VPWR _01414_ sky130_fd_sc_hd__mux2_1
XFILLER_27_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06874_ data_array.data0\[12\]\[12\] net1388 net1294 data_array.data0\[15\]\[12\]
+ _04166_ VGND VGND VPWR VPWR _04167_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_2_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08613_ net773 net4125 net523 VGND VGND VPWR VPWR _00372_ sky130_fd_sc_hd__mux2_1
X_05825_ _03247_ _03288_ VGND VGND VPWR VPWR _03342_ sky130_fd_sc_hd__or2_1
X_09593_ net977 net4133 net399 VGND VGND VPWR VPWR _01345_ sky130_fd_sc_hd__mux2_1
X_08544_ net779 net4034 net582 VGND VGND VPWR VPWR _00312_ sky130_fd_sc_hd__mux2_1
XFILLER_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05756_ fsm.tag_out1\[10\] net9 VGND VGND VPWR VPWR _03273_ sky130_fd_sc_hd__and2b_1
XFILLER_24_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08475_ net824 _05552_ VGND VGND VPWR VPWR _05553_ sky130_fd_sc_hd__or2_1
XFILLER_165_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05687_ net17 fsm.tag_out0\[17\] VGND VGND VPWR VPWR _03204_ sky130_fd_sc_hd__and2b_1
XFILLER_39_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07426_ data_array.data0\[0\]\[62\] net1412 net1318 data_array.data0\[3\]\[62\] _04668_
+ VGND VGND VPWR VPWR _04669_ sky130_fd_sc_hd__a221o_1
XFILLER_51_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07357_ data_array.data0\[9\]\[56\] net1531 net1435 data_array.data0\[10\]\[56\]
+ VGND VGND VPWR VPWR _04606_ sky130_fd_sc_hd__a22o_1
XFILLER_148_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06308_ tag_array.tag0\[13\]\[11\] net1593 net1497 tag_array.tag0\[14\]\[11\] VGND
+ VGND VPWR VPWR _03652_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_21_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07288_ data_array.data0\[8\]\[50\] net1346 net1252 data_array.data0\[11\]\[50\]
+ _04542_ VGND VGND VPWR VPWR _04543_ sky130_fd_sc_hd__a221o_1
XFILLER_164_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09027_ net2024 net917 net422 VGND VGND VPWR VPWR _00782_ sky130_fd_sc_hd__mux2_1
X_06239_ net1626 _03583_ _03587_ net1200 VGND VGND VPWR VPWR _03590_ sky130_fd_sc_hd__a22o_1
XFILLER_105_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_938 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold250 data_array.data1\[4\]\[22\] VGND VGND VPWR VPWR net1901 sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 data_array.data0\[4\]\[6\] VGND VGND VPWR VPWR net1912 sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 tag_array.tag1\[4\]\[0\] VGND VGND VPWR VPWR net1923 sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 tag_array.tag1\[0\]\[21\] VGND VGND VPWR VPWR net1934 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 data_array.data0\[8\]\[57\] VGND VGND VPWR VPWR net1945 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout730 _05395_ VGND VGND VPWR VPWR net730 sky130_fd_sc_hd__clkbuf_2
Xfanout741 _05391_ VGND VGND VPWR VPWR net741 sky130_fd_sc_hd__buf_1
XFILLER_104_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09929_ net807 _05583_ VGND VGND VPWR VPWR _03127_ sky130_fd_sc_hd__nand2_8
Xfanout752 net753 VGND VGND VPWR VPWR net752 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_130_Right_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout763 _05379_ VGND VGND VPWR VPWR net763 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_146_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout774 net775 VGND VGND VPWR VPWR net774 sky130_fd_sc_hd__clkbuf_2
Xfanout785 _05369_ VGND VGND VPWR VPWR net785 sky130_fd_sc_hd__buf_1
Xfanout796 net797 VGND VGND VPWR VPWR net796 sky130_fd_sc_hd__clkbuf_8
X_12940_ clknet_leaf_84_clk _01634_ VGND VGND VPWR VPWR data_array.data0\[13\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_107_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ clknet_leaf_234_clk _01565_ VGND VGND VPWR VPWR data_array.data0\[12\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_142_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ clknet_leaf_92_clk _00630_ VGND VGND VPWR VPWR data_array.data0\[7\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_103_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11753_ clknet_leaf_60_clk _00561_ VGND VGND VPWR VPWR data_array.data0\[8\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ net2811 net900 net481 VGND VGND VPWR VPWR _02449_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_120_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14472_ clknet_leaf_9_clk _03095_ VGND VGND VPWR VPWR data_array.data1\[7\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
X_11684_ clknet_leaf_96_clk _00492_ VGND VGND VPWR VPWR tag_array.tag1\[15\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_10635_ net2045 net922 net473 VGND VGND VPWR VPWR _02380_ sky130_fd_sc_hd__mux2_1
X_13423_ clknet_leaf_44_clk _02053_ VGND VGND VPWR VPWR data_array.data1\[8\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_139_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload109 clknet_leaf_92_clk VGND VGND VPWR VPWR clkload109/Y sky130_fd_sc_hd__clkinvlp_4
X_13354_ clknet_leaf_224_clk _01984_ VGND VGND VPWR VPWR data_array.data0\[10\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
X_10566_ net943 net4513 net462 VGND VGND VPWR VPWR _02311_ sky130_fd_sc_hd__mux2_1
XFILLER_127_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12305_ clknet_leaf_166_clk _01063_ VGND VGND VPWR VPWR tag_array.tag1\[12\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_182_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13285_ clknet_leaf_207_clk _01915_ VGND VGND VPWR VPWR data_array.data0\[11\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_127_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10497_ net957 net3375 net349 VGND VGND VPWR VPWR _02242_ sky130_fd_sc_hd__mux2_1
XFILLER_182_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12236_ clknet_leaf_150_clk _00165_ VGND VGND VPWR VPWR fsm.tag_out1\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_166_3545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_166_3556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12167_ clknet_leaf_182_clk _00975_ VGND VGND VPWR VPWR tag_array.tag0\[13\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11118_ net1045 net4018 net545 VGND VGND VPWR VPWR _02861_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_183_3870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_3881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12098_ clknet_leaf_78_clk _00906_ VGND VGND VPWR VPWR data_array.data1\[14\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_127_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11049_ net2763 net1064 net334 VGND VGND VPWR VPWR _02792_ sky130_fd_sc_hd__mux2_1
Xinput7 cpu_addr[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_2
XFILLER_76_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06590_ tag_array.tag1\[0\]\[11\] net1385 net1291 tag_array.tag1\[3\]\[11\] _03908_
+ VGND VGND VPWR VPWR _03909_ sky130_fd_sc_hd__a221o_1
XFILLER_64_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08260_ net1649 net1160 net22 VGND VGND VPWR VPWR _05408_ sky130_fd_sc_hd__and3_1
XFILLER_33_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07211_ data_array.data0\[8\]\[43\] net1377 net1283 data_array.data0\[11\]\[43\]
+ _04472_ VGND VGND VPWR VPWR _04473_ sky130_fd_sc_hd__a221o_1
X_08191_ net1279 net1172 VGND VGND VPWR VPWR _05361_ sky130_fd_sc_hd__nand2_1
XFILLER_158_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07142_ net1183 _04405_ _04409_ net1231 VGND VGND VPWR VPWR _04411_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_41_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07073_ data_array.data0\[1\]\[30\] net1581 net1485 data_array.data0\[2\]\[30\] VGND
+ VGND VPWR VPWR _04348_ sky130_fd_sc_hd__a22o_1
XFILLER_106_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput300 net300 VGND VGND VPWR VPWR mem_wdata[43] sky130_fd_sc_hd__buf_2
Xoutput311 net311 VGND VGND VPWR VPWR mem_wdata[53] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_144_Left_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput322 net322 VGND VGND VPWR VPWR mem_wdata[63] sky130_fd_sc_hd__buf_2
X_06024_ net1162 net12 VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__and2_1
XFILLER_133_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07975_ data_array.data1\[1\]\[48\] net1583 net1487 data_array.data1\[2\]\[48\] VGND
+ VGND VPWR VPWR _05168_ sky130_fd_sc_hd__a22o_1
XFILLER_102_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06926_ data_array.data0\[1\]\[17\] net1530 net1434 data_array.data0\[2\]\[17\] VGND
+ VGND VPWR VPWR _04214_ sky130_fd_sc_hd__a22o_1
X_09714_ net732 net2935 net610 VGND VGND VPWR VPWR _01466_ sky130_fd_sc_hd__mux2_1
XFILLER_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09645_ net709 net2069 net616 VGND VGND VPWR VPWR _01397_ sky130_fd_sc_hd__mux2_1
X_06857_ _04150_ _04151_ VGND VGND VPWR VPWR _00001_ sky130_fd_sc_hd__or2_1
XFILLER_16_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_153_Left_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_915 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05808_ _03169_ _03185_ _03208_ _03224_ VGND VGND VPWR VPWR _03325_ sky130_fd_sc_hd__or4_1
X_09576_ net1046 net3842 net397 VGND VGND VPWR VPWR _01328_ sky130_fd_sc_hd__mux2_1
XFILLER_71_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06788_ data_array.data0\[0\]\[4\] net1391 net1297 data_array.data0\[3\]\[4\] _04088_
+ VGND VGND VPWR VPWR _04089_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_65_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08527_ net1719 net593 VGND VGND VPWR VPWR _00303_ sky130_fd_sc_hd__nand2b_1
X_05739_ net5 _03138_ net15 _03141_ VGND VGND VPWR VPWR _03256_ sky130_fd_sc_hd__a22o_1
Xclkbuf_5_20__f_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_5_20__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_24_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08458_ net1126 _05541_ VGND VGND VPWR VPWR _05542_ sky130_fd_sc_hd__and2_2
X_07409_ data_array.data0\[12\]\[61\] net1361 net1267 data_array.data0\[15\]\[61\]
+ _04652_ VGND VGND VPWR VPWR _04653_ sky130_fd_sc_hd__a221o_1
X_08389_ net1127 _05495_ VGND VGND VPWR VPWR _05496_ sky130_fd_sc_hd__and2_1
XFILLER_183_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10420_ net1859 net974 net663 VGND VGND VPWR VPWR _02166_ sky130_fd_sc_hd__mux2_1
XFILLER_137_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_162_Left_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10351_ net694 net3472 net591 VGND VGND VPWR VPWR _02098_ sky130_fd_sc_hd__mux2_1
XFILLER_136_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13070_ clknet_leaf_221_clk _01764_ VGND VGND VPWR VPWR data_array.data1\[13\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_10282_ net2661 net1034 net640 VGND VGND VPWR VPWR _02029_ sky130_fd_sc_hd__mux2_1
XFILLER_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12021_ clknet_leaf_34_clk _00829_ VGND VGND VPWR VPWR data_array.data0\[6\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_116_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1503 net1504 VGND VGND VPWR VPWR net1503 sky130_fd_sc_hd__buf_2
Xfanout1514 net1516 VGND VGND VPWR VPWR net1514 sky130_fd_sc_hd__clkbuf_4
Xfanout1525 net1526 VGND VGND VPWR VPWR net1525 sky130_fd_sc_hd__clkbuf_4
Xfanout1536 net1543 VGND VGND VPWR VPWR net1536 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_144_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1547 net1549 VGND VGND VPWR VPWR net1547 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_144_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout560 _05593_ VGND VGND VPWR VPWR net560 sky130_fd_sc_hd__clkbuf_4
Xfanout1558 net1560 VGND VGND VPWR VPWR net1558 sky130_fd_sc_hd__clkbuf_4
Xfanout571 net572 VGND VGND VPWR VPWR net571 sky130_fd_sc_hd__buf_4
Xfanout1569 net1573 VGND VGND VPWR VPWR net1569 sky130_fd_sc_hd__clkbuf_2
Xfanout582 net584 VGND VGND VPWR VPWR net582 sky130_fd_sc_hd__clkbuf_8
XFILLER_65_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_161_3453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout593 net594 VGND VGND VPWR VPWR net593 sky130_fd_sc_hd__buf_2
X_13972_ clknet_leaf_86_clk _02601_ VGND VGND VPWR VPWR data_array.data1\[5\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_161_3464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_171_Left_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12923_ clknet_leaf_237_clk _01617_ VGND VGND VPWR VPWR data_array.data0\[13\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_73_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12854_ clknet_leaf_22_clk _01548_ VGND VGND VPWR VPWR data_array.data0\[12\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11805_ clknet_leaf_112_clk _00613_ VGND VGND VPWR VPWR data_array.data0\[7\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_12785_ clknet_leaf_191_clk _01479_ VGND VGND VPWR VPWR tag_array.tag1\[10\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_92_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11736_ clknet_leaf_248_clk _00544_ VGND VGND VPWR VPWR data_array.data0\[8\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_25_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14455_ clknet_leaf_240_clk _03078_ VGND VGND VPWR VPWR data_array.data1\[7\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
X_11667_ clknet_leaf_139_clk _00475_ VGND VGND VPWR VPWR tag_array.tag1\[1\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_180_Left_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13406_ clknet_leaf_250_clk _02036_ VGND VGND VPWR VPWR data_array.data1\[8\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10618_ net1974 net990 net472 VGND VGND VPWR VPWR _02363_ sky130_fd_sc_hd__mux2_1
X_14386_ clknet_leaf_118_clk _03009_ VGND VGND VPWR VPWR data_array.data1\[10\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
X_11598_ clknet_leaf_167_clk _00406_ VGND VGND VPWR VPWR tag_array.tag1\[4\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_10549_ net1010 net3970 net453 VGND VGND VPWR VPWR _02294_ sky130_fd_sc_hd__mux2_1
X_13337_ clknet_leaf_23_clk _01967_ VGND VGND VPWR VPWR data_array.data0\[10\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13268_ clknet_leaf_259_clk _01898_ VGND VGND VPWR VPWR data_array.data0\[11\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_69_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12219_ clknet_leaf_151_clk _00167_ VGND VGND VPWR VPWR fsm.tag_out1\[1\] sky130_fd_sc_hd__dfxtp_1
X_13199_ clknet_leaf_118_clk _00093_ VGND VGND VPWR VPWR data_array.rdata1\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_37_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2409 tag_array.tag1\[13\]\[3\] VGND VGND VPWR VPWR net4060 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_181_3829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1708 tag_array.tag0\[8\]\[22\] VGND VGND VPWR VPWR net3359 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1719 tag_array.tag1\[12\]\[13\] VGND VGND VPWR VPWR net3370 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07760_ data_array.data1\[13\]\[29\] net1577 net1481 data_array.data1\[14\]\[29\]
+ VGND VGND VPWR VPWR _04972_ sky130_fd_sc_hd__a22o_1
XFILLER_96_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06711_ tag_array.tag1\[4\]\[22\] net1362 net1268 tag_array.tag1\[7\]\[22\] _04018_
+ VGND VGND VPWR VPWR _04019_ sky130_fd_sc_hd__a221o_1
X_07691_ net1619 _04903_ _04907_ net1193 VGND VGND VPWR VPWR _04910_ sky130_fd_sc_hd__a22o_1
XFILLER_38_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09430_ net945 net3673 net578 VGND VGND VPWR VPWR _01183_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_200_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_200_clk
+ sky130_fd_sc_hd__clkbuf_8
X_06642_ tag_array.tag1\[9\]\[16\] net1608 net1512 tag_array.tag1\[10\]\[16\] VGND
+ VGND VPWR VPWR _03956_ sky130_fd_sc_hd__a22o_1
XFILLER_24_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09361_ net956 net4559 net406 VGND VGND VPWR VPWR _01114_ sky130_fd_sc_hd__mux2_1
XFILLER_24_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06573_ tag_array.tag1\[12\]\[10\] net1404 net1310 tag_array.tag1\[15\]\[10\] _03892_
+ VGND VGND VPWR VPWR _03893_ sky130_fd_sc_hd__a221o_1
XFILLER_80_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_970 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08312_ net1906 net1060 net693 VGND VGND VPWR VPWR _00233_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09292_ net710 net4402 net556 VGND VGND VPWR VPWR _01046_ sky130_fd_sc_hd__mux2_1
XFILLER_166_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_12 _03127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_23 _03515_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08243_ fsm.tag_out1\[16\] net817 net809 fsm.tag_out0\[16\] _05396_ VGND VGND VPWR
+ VPWR _05397_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_60_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_34 net381 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_45 net594 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_56 net1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_67 net1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08174_ lru_array.lru_mem\[0\] net1371 net1277 lru_array.lru_mem\[3\] _05348_ VGND
+ VGND VPWR VPWR _05349_ sky130_fd_sc_hd__a221o_1
XANTENNA_78 net417 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_89 net1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_267_clk clknet_5_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_267_clk
+ sky130_fd_sc_hd__clkbuf_8
X_07125_ data_array.data0\[4\]\[35\] net1346 net1252 data_array.data0\[7\]\[35\] _04394_
+ VGND VGND VPWR VPWR _04395_ sky130_fd_sc_hd__a221o_1
XFILLER_118_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07056_ data_array.data0\[13\]\[29\] net1571 net1475 data_array.data0\[14\]\[29\]
+ VGND VGND VPWR VPWR _04332_ sky130_fd_sc_hd__a22o_1
XFILLER_134_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06007_ net152 net1152 _03464_ _03465_ VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__a22o_1
XFILLER_115_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput174 net174 VGND VGND VPWR VPWR cpu_rdata[18] sky130_fd_sc_hd__buf_2
XFILLER_0_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput185 net185 VGND VGND VPWR VPWR cpu_rdata[28] sky130_fd_sc_hd__buf_2
Xoutput196 net196 VGND VGND VPWR VPWR cpu_rdata[38] sky130_fd_sc_hd__buf_6
Xhold2910 data_array.data1\[6\]\[21\] VGND VGND VPWR VPWR net4561 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2921 data_array.data1\[11\]\[38\] VGND VGND VPWR VPWR net4572 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2932 data_array.data1\[15\]\[28\] VGND VGND VPWR VPWR net4583 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2943 data_array.data1\[11\]\[22\] VGND VGND VPWR VPWR net4594 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2954 data_array.data1\[3\]\[28\] VGND VGND VPWR VPWR net4605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2965 tag_array.tag1\[10\]\[1\] VGND VGND VPWR VPWR net4616 sky130_fd_sc_hd__dlygate4sd3_1
X_07958_ data_array.data1\[9\]\[47\] net1589 net1493 data_array.data1\[10\]\[47\]
+ VGND VGND VPWR VPWR _05152_ sky130_fd_sc_hd__a22o_1
XFILLER_102_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06909_ data_array.data0\[0\]\[15\] net1390 net1296 data_array.data0\[3\]\[15\] _04198_
+ VGND VGND VPWR VPWR _04199_ sky130_fd_sc_hd__a221o_1
XFILLER_56_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07889_ net1209 _05083_ _05087_ net1635 VGND VGND VPWR VPWR _05090_ sky130_fd_sc_hd__a22o_1
XFILLER_46_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09628_ net776 net2967 net615 VGND VGND VPWR VPWR _01380_ sky130_fd_sc_hd__mux2_1
X_09559_ _05414_ _05595_ VGND VGND VPWR VPWR _03124_ sky130_fd_sc_hd__or2_1
XFILLER_102_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12570_ clknet_leaf_170_clk _01264_ VGND VGND VPWR VPWR tag_array.tag0\[10\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11521_ clknet_leaf_231_clk _00329_ VGND VGND VPWR VPWR tag_array.tag1\[9\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11452_ clknet_leaf_260_clk _00262_ VGND VGND VPWR VPWR data_array.data0\[0\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
X_14240_ clknet_leaf_87_clk _02869_ VGND VGND VPWR VPWR data_array.data1\[12\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_258_clk clknet_5_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_258_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10403_ net1785 net1040 net661 VGND VGND VPWR VPWR _02149_ sky130_fd_sc_hd__mux2_1
X_14171_ clknet_leaf_60_clk _02800_ VGND VGND VPWR VPWR data_array.data0\[2\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_11383_ net164 VGND VGND VPWR VPWR _00193_ sky130_fd_sc_hd__inv_2
XFILLER_109_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_78_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13122_ clknet_leaf_160_clk _01816_ VGND VGND VPWR VPWR tag_array.tag0\[3\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_10334_ net763 net4337 net592 VGND VGND VPWR VPWR _02081_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_115_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13053_ clknet_leaf_68_clk _01747_ VGND VGND VPWR VPWR data_array.data1\[13\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_10265_ net2708 net1101 net634 VGND VGND VPWR VPWR _02012_ sky130_fd_sc_hd__mux2_1
XFILLER_3_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_163_3504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1300 net1306 VGND VGND VPWR VPWR net1300 sky130_fd_sc_hd__clkbuf_4
XFILLER_87_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12004_ clknet_leaf_49_clk _00812_ VGND VGND VPWR VPWR data_array.data0\[6\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_121_931 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1311 net1312 VGND VGND VPWR VPWR net1311 sky130_fd_sc_hd__clkbuf_4
XFILLER_87_75 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1322 net1328 VGND VGND VPWR VPWR net1322 sky130_fd_sc_hd__buf_2
X_10196_ net1023 net3601 net355 VGND VGND VPWR VPWR _01943_ sky130_fd_sc_hd__mux2_1
XFILLER_78_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1333 net1334 VGND VGND VPWR VPWR net1333 sky130_fd_sc_hd__clkbuf_4
Xfanout1344 net1345 VGND VGND VPWR VPWR net1344 sky130_fd_sc_hd__clkbuf_4
Xfanout1355 net1364 VGND VGND VPWR VPWR net1355 sky130_fd_sc_hd__buf_2
XFILLER_66_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1001 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1366 net1367 VGND VGND VPWR VPWR net1366 sky130_fd_sc_hd__clkbuf_4
XFILLER_121_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1377 net1378 VGND VGND VPWR VPWR net1377 sky130_fd_sc_hd__clkbuf_4
Xfanout390 net392 VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__clkbuf_8
Xfanout1388 net1400 VGND VGND VPWR VPWR net1388 sky130_fd_sc_hd__clkbuf_4
Xfanout1399 net1400 VGND VGND VPWR VPWR net1399 sky130_fd_sc_hd__clkbuf_4
XFILLER_98_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13955_ clknet_leaf_55_clk _02584_ VGND VGND VPWR VPWR data_array.data1\[4\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
X_12906_ clknet_leaf_111_clk _01600_ VGND VGND VPWR VPWR data_array.data0\[13\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_13886_ clknet_leaf_214_clk _02515_ VGND VGND VPWR VPWR data_array.data1\[3\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12837_ clknet_leaf_203_clk _01531_ VGND VGND VPWR VPWR data_array.data0\[12\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_178_3780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12768_ clknet_leaf_166_clk _01462_ VGND VGND VPWR VPWR tag_array.tag0\[6\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_175_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11719_ clknet_leaf_107_clk _00527_ VGND VGND VPWR VPWR tag_array.tag0\[9\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_175_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_174_3699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12699_ clknet_leaf_108_clk _01393_ VGND VGND VPWR VPWR tag_array.tag0\[8\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_14438_ clknet_leaf_24_clk _03061_ VGND VGND VPWR VPWR data_array.data1\[7\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput10 cpu_addr[18] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_2
Xinput21 cpu_addr[28] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput32 cpu_addr[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_2
Xinput43 cpu_wdata[18] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_249_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_249_clk
+ sky130_fd_sc_hd__clkbuf_8
Xinput54 cpu_wdata[28] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_1
Xinput65 cpu_wdata[38] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_1
X_14369_ clknet_leaf_67_clk _02992_ VGND VGND VPWR VPWR data_array.data1\[10\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold805 tag_array.tag1\[10\]\[10\] VGND VGND VPWR VPWR net2456 sky130_fd_sc_hd__dlygate4sd3_1
Xinput76 cpu_wdata[48] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__clkbuf_1
Xhold816 tag_array.tag0\[6\]\[20\] VGND VGND VPWR VPWR net2467 sky130_fd_sc_hd__dlygate4sd3_1
Xinput87 cpu_wdata[58] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_1
XFILLER_155_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput98 cpu_write VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__buf_4
Xhold827 data_array.data1\[9\]\[14\] VGND VGND VPWR VPWR net2478 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold838 data_array.data0\[14\]\[49\] VGND VGND VPWR VPWR net2489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold849 data_array.data0\[1\]\[58\] VGND VGND VPWR VPWR net2500 sky130_fd_sc_hd__dlygate4sd3_1
X_08930_ net1047 net4074 net428 VGND VGND VPWR VPWR _00686_ sky130_fd_sc_hd__mux2_1
XFILLER_112_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2206 data_array.data1\[11\]\[17\] VGND VGND VPWR VPWR net3857 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2217 data_array.data0\[11\]\[45\] VGND VGND VPWR VPWR net3868 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2228 tag_array.tag0\[11\]\[6\] VGND VGND VPWR VPWR net3879 sky130_fd_sc_hd__dlygate4sd3_1
X_08861_ net1060 net3896 net440 VGND VGND VPWR VPWR _00618_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2239 data_array.data0\[6\]\[42\] VGND VGND VPWR VPWR net3890 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1505 tag_array.tag0\[2\]\[16\] VGND VGND VPWR VPWR net3156 sky130_fd_sc_hd__dlygate4sd3_1
X_07812_ net1206 _05013_ _05017_ net1632 VGND VGND VPWR VPWR _05020_ sky130_fd_sc_hd__a22o_1
Xhold1516 data_array.data1\[7\]\[41\] VGND VGND VPWR VPWR net3167 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1527 data_array.data1\[12\]\[26\] VGND VGND VPWR VPWR net3178 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08792_ net1878 net1076 net443 VGND VGND VPWR VPWR _00550_ sky130_fd_sc_hd__mux2_1
XFILLER_69_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1538 tag_array.tag0\[14\]\[16\] VGND VGND VPWR VPWR net3189 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1549 data_array.data0\[13\]\[26\] VGND VGND VPWR VPWR net3200 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_42_1062 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07743_ data_array.data1\[12\]\[27\] net1358 net1264 data_array.data1\[15\]\[27\]
+ _04956_ VGND VGND VPWR VPWR _04957_ sky130_fd_sc_hd__a221o_1
XFILLER_38_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07674_ data_array.data1\[1\]\[21\] net1555 net1459 data_array.data1\[2\]\[21\] VGND
+ VGND VPWR VPWR _04894_ sky130_fd_sc_hd__a22o_1
XFILLER_53_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06625_ net1222 _03935_ _03939_ net1173 VGND VGND VPWR VPWR _03941_ sky130_fd_sc_hd__a22o_1
X_09413_ net1014 net3725 net586 VGND VGND VPWR VPWR _01166_ sky130_fd_sc_hd__mux2_1
XFILLER_53_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06556_ tag_array.tag1\[1\]\[8\] net1608 net1512 tag_array.tag1\[2\]\[8\] VGND VGND
+ VPWR VPWR _03878_ sky130_fd_sc_hd__a22o_1
X_09344_ net1026 net4196 net404 VGND VGND VPWR VPWR _01097_ sky130_fd_sc_hd__mux2_1
XFILLER_178_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09275_ net778 net4060 net559 VGND VGND VPWR VPWR _01029_ sky130_fd_sc_hd__mux2_1
X_06487_ tag_array.tag1\[4\]\[2\] net1351 net1257 tag_array.tag1\[7\]\[2\] _03814_
+ VGND VGND VPWR VPWR _03815_ sky130_fd_sc_hd__a221o_1
XFILLER_20_163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08226_ net750 net3293 net805 VGND VGND VPWR VPWR _00206_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_99_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08157_ tag_array.dirty0\[12\] net1403 net1309 tag_array.dirty0\[15\] _05332_ VGND
+ VGND VPWR VPWR _05333_ sky130_fd_sc_hd__a221o_1
XFILLER_113_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07108_ net1205 _04373_ _04377_ net1631 VGND VGND VPWR VPWR _04380_ sky130_fd_sc_hd__a22o_1
X_08088_ net1171 _05265_ _05269_ net1219 VGND VGND VPWR VPWR _05271_ sky130_fd_sc_hd__a22o_1
XFILLER_162_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07039_ data_array.data0\[12\]\[27\] net1347 net1253 data_array.data0\[15\]\[27\]
+ _04316_ VGND VGND VPWR VPWR _04317_ sky130_fd_sc_hd__a221o_1
X_10050_ net887 net3497 net556 VGND VGND VPWR VPWR _01799_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_73_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_110_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2740 data_array.data1\[11\]\[47\] VGND VGND VPWR VPWR net4391 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2751 tag_array.tag1\[13\]\[20\] VGND VGND VPWR VPWR net4402 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2762 tag_array.tag1\[3\]\[9\] VGND VGND VPWR VPWR net4413 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2773 data_array.data0\[6\]\[27\] VGND VGND VPWR VPWR net4424 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2784 tag_array.tag0\[8\]\[8\] VGND VGND VPWR VPWR net4435 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2795 data_array.data0\[15\]\[14\] VGND VGND VPWR VPWR net4446 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13740_ clknet_leaf_83_clk _02369_ VGND VGND VPWR VPWR data_array.data1\[1\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_27_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10952_ net934 net3628 net533 VGND VGND VPWR VPWR _02697_ sky130_fd_sc_hd__mux2_1
XFILLER_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13671_ clknet_leaf_37_clk _02300_ VGND VGND VPWR VPWR data_array.data1\[15\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_10883_ net953 net3594 net515 VGND VGND VPWR VPWR _02628_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_139_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12622_ clknet_leaf_71_clk _01316_ VGND VGND VPWR VPWR data_array.data0\[15\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_58_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_156_3363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12553_ clknet_leaf_107_clk _01247_ VGND VGND VPWR VPWR tag_array.tag0\[11\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_169_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_664 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11504_ clknet_leaf_191_clk _00312_ VGND VGND VPWR VPWR tag_array.tag1\[9\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12484_ clknet_leaf_118_clk _01178_ VGND VGND VPWR VPWR data_array.data1\[9\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14223_ clknet_leaf_118_clk _02852_ VGND VGND VPWR VPWR data_array.data1\[12\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11435_ clknet_leaf_92_clk _00245_ VGND VGND VPWR VPWR data_array.data0\[0\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14154_ clknet_leaf_247_clk _02783_ VGND VGND VPWR VPWR data_array.data0\[2\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_11366_ net1646 net3525 net606 VGND VGND VPWR VPWR _03109_ sky130_fd_sc_hd__mux2_1
XFILLER_180_661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10317_ net2175 net893 net634 VGND VGND VPWR VPWR _02064_ sky130_fd_sc_hd__mux2_1
X_13105_ clknet_leaf_21_clk _01799_ VGND VGND VPWR VPWR data_array.data1\[13\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_130_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11297_ net1104 net4292 net795 VGND VGND VPWR VPWR _03040_ sky130_fd_sc_hd__mux2_1
X_14085_ clknet_leaf_211_clk _02714_ VGND VGND VPWR VPWR data_array.data1\[6\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_152_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13036_ clknet_leaf_1_clk _01730_ VGND VGND VPWR VPWR data_array.data0\[3\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
X_10248_ net751 net3973 net596 VGND VGND VPWR VPWR _01995_ sky130_fd_sc_hd__mux2_1
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1130 _05418_ VGND VGND VPWR VPWR net1130 sky130_fd_sc_hd__buf_6
XFILLER_66_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1141 _03477_ VGND VGND VPWR VPWR net1141 sky130_fd_sc_hd__clkbuf_8
XFILLER_113_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10179_ net1088 net2185 net356 VGND VGND VPWR VPWR _01926_ sky130_fd_sc_hd__mux2_1
Xfanout1152 net1153 VGND VGND VPWR VPWR net1152 sky130_fd_sc_hd__clkbuf_4
XFILLER_26_1079 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1163 net1164 VGND VGND VPWR VPWR net1163 sky130_fd_sc_hd__clkbuf_2
Xfanout1174 net1175 VGND VGND VPWR VPWR net1174 sky130_fd_sc_hd__buf_4
Xfanout1185 net1186 VGND VGND VPWR VPWR net1185 sky130_fd_sc_hd__clkbuf_2
Xfanout1196 net1198 VGND VGND VPWR VPWR net1196 sky130_fd_sc_hd__buf_4
XFILLER_47_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13938_ clknet_leaf_87_clk _02567_ VGND VGND VPWR VPWR data_array.data1\[4\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_176_3739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13869_ clknet_leaf_214_clk _02498_ VGND VGND VPWR VPWR data_array.data1\[3\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
X_06410_ tag_array.tag0\[4\]\[20\] net1369 net1275 tag_array.tag0\[7\]\[20\] _03744_
+ VGND VGND VPWR VPWR _03745_ sky130_fd_sc_hd__a221o_1
XFILLER_50_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07390_ data_array.data0\[13\]\[59\] net1570 net1474 data_array.data0\[14\]\[59\]
+ VGND VGND VPWR VPWR _04636_ sky130_fd_sc_hd__a22o_1
X_06341_ tag_array.tag0\[9\]\[14\] net1559 net1463 tag_array.tag0\[10\]\[14\] VGND
+ VGND VPWR VPWR _03682_ sky130_fd_sc_hd__a22o_1
XFILLER_176_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_962 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09060_ net1047 net2681 net412 VGND VGND VPWR VPWR _00814_ sky130_fd_sc_hd__mux2_1
X_06272_ net1634 _03613_ _03617_ net1208 VGND VGND VPWR VPWR _03620_ sky130_fd_sc_hd__a22o_1
X_08011_ net1167 _05195_ _05199_ net1215 VGND VGND VPWR VPWR _05201_ sky130_fd_sc_hd__a22o_1
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold602 data_array.data1\[1\]\[34\] VGND VGND VPWR VPWR net2253 sky130_fd_sc_hd__dlygate4sd3_1
Xhold613 data_array.data0\[8\]\[36\] VGND VGND VPWR VPWR net2264 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold624 data_array.data0\[4\]\[23\] VGND VGND VPWR VPWR net2275 sky130_fd_sc_hd__dlygate4sd3_1
Xhold635 data_array.data0\[5\]\[15\] VGND VGND VPWR VPWR net2286 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold646 data_array.data0\[0\]\[45\] VGND VGND VPWR VPWR net2297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 tag_array.tag0\[2\]\[24\] VGND VGND VPWR VPWR net2308 sky130_fd_sc_hd__dlygate4sd3_1
Xhold668 data_array.data1\[0\]\[42\] VGND VGND VPWR VPWR net2319 sky130_fd_sc_hd__dlygate4sd3_1
X_09962_ net983 net3908 net370 VGND VGND VPWR VPWR _01711_ sky130_fd_sc_hd__mux2_1
XFILLER_131_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold679 tag_array.tag1\[2\]\[8\] VGND VGND VPWR VPWR net2330 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2003 data_array.data0\[15\]\[54\] VGND VGND VPWR VPWR net3654 sky130_fd_sc_hd__dlygate4sd3_1
X_08913_ net807 _05577_ VGND VGND VPWR VPWR _05609_ sky130_fd_sc_hd__nand2_1
X_09893_ net897 net4433 net378 VGND VGND VPWR VPWR _01643_ sky130_fd_sc_hd__mux2_1
XFILLER_69_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2014 tag_array.tag0\[14\]\[12\] VGND VGND VPWR VPWR net3665 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2025 tag_array.tag0\[10\]\[11\] VGND VGND VPWR VPWR net3676 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2036 data_array.data0\[12\]\[8\] VGND VGND VPWR VPWR net3687 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1302 tag_array.tag1\[3\]\[5\] VGND VGND VPWR VPWR net2953 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2047 data_array.data0\[15\]\[47\] VGND VGND VPWR VPWR net3698 sky130_fd_sc_hd__dlygate4sd3_1
X_08844_ net1978 net869 net449 VGND VGND VPWR VPWR _00602_ sky130_fd_sc_hd__mux2_1
Xhold1313 data_array.data0\[8\]\[33\] VGND VGND VPWR VPWR net2964 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2058 data_array.data1\[9\]\[4\] VGND VGND VPWR VPWR net3709 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2069 tag_array.tag0\[8\]\[19\] VGND VGND VPWR VPWR net3720 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1324 tag_array.tag0\[12\]\[19\] VGND VGND VPWR VPWR net2975 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1335 data_array.data0\[12\]\[25\] VGND VGND VPWR VPWR net2986 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1346 data_array.data1\[1\]\[37\] VGND VGND VPWR VPWR net2997 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1357 data_array.data1\[5\]\[41\] VGND VGND VPWR VPWR net3008 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05987_ data_array.rdata0\[52\] net848 net1144 VGND VGND VPWR VPWR _03452_ sky130_fd_sc_hd__o21a_1
XFILLER_84_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1368 data_array.data1\[5\]\[24\] VGND VGND VPWR VPWR net3019 sky130_fd_sc_hd__dlygate4sd3_1
X_08775_ net722 net4007 net451 VGND VGND VPWR VPWR _00534_ sky130_fd_sc_hd__mux2_1
XFILLER_26_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1379 data_array.data1\[2\]\[21\] VGND VGND VPWR VPWR net3030 sky130_fd_sc_hd__dlygate4sd3_1
X_07726_ _04940_ _04941_ VGND VGND VPWR VPWR _00081_ sky130_fd_sc_hd__or2_1
X_07657_ data_array.data1\[0\]\[19\] net1394 net1300 data_array.data1\[3\]\[19\] _04878_
+ VGND VGND VPWR VPWR _04879_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_0_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06608_ tag_array.tag1\[4\]\[13\] net1420 net1326 tag_array.tag1\[7\]\[13\] _03924_
+ VGND VGND VPWR VPWR _03925_ sky130_fd_sc_hd__a221o_1
XFILLER_13_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07588_ data_array.data1\[9\]\[13\] net1551 net1455 data_array.data1\[10\]\[13\]
+ VGND VGND VPWR VPWR _04816_ sky130_fd_sc_hd__a22o_1
XFILLER_43_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06539_ tag_array.tag1\[9\]\[7\] net1611 net1515 tag_array.tag1\[10\]\[7\] VGND VGND
+ VPWR VPWR _03862_ sky130_fd_sc_hd__a22o_1
X_09327_ net1093 net3783 net407 VGND VGND VPWR VPWR _01080_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09258_ net746 net4387 net575 VGND VGND VPWR VPWR _01012_ sky130_fd_sc_hd__mux2_1
XFILLER_154_606 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08209_ net1650 net1163 net4 VGND VGND VPWR VPWR _05374_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_151_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09189_ net723 net4469 net628 VGND VGND VPWR VPWR _00943_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_151_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_177_Right_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11220_ net893 net3103 net649 VGND VGND VPWR VPWR _02963_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11151_ net915 net2825 net549 VGND VGND VPWR VPWR _02894_ sky130_fd_sc_hd__mux2_1
XFILLER_175_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10102_ net3080 net715 net639 VGND VGND VPWR VPWR _01851_ sky130_fd_sc_hd__mux2_1
XFILLER_122_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11082_ net2656 net932 _03133_ VGND VGND VPWR VPWR _02825_ sky130_fd_sc_hd__mux2_1
XFILLER_68_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10033_ net953 net4611 net557 VGND VGND VPWR VPWR _01782_ sky130_fd_sc_hd__mux2_1
XFILLER_76_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2570 tag_array.tag1\[3\]\[13\] VGND VGND VPWR VPWR net4221 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2581 data_array.data0\[10\]\[16\] VGND VGND VPWR VPWR net4232 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_64_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2592 tag_array.tag0\[12\]\[7\] VGND VGND VPWR VPWR net4243 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_64_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1880 data_array.data1\[9\]\[49\] VGND VGND VPWR VPWR net3531 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1891 data_array.data1\[9\]\[31\] VGND VGND VPWR VPWR net3542 sky130_fd_sc_hd__dlygate4sd3_1
X_11984_ clknet_leaf_209_clk _00792_ VGND VGND VPWR VPWR data_array.data0\[4\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_158_3403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13723_ clknet_leaf_66_clk _02352_ VGND VGND VPWR VPWR data_array.data1\[1\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_10935_ net1000 net3258 net528 VGND VGND VPWR VPWR _02680_ sky130_fd_sc_hd__mux2_1
XFILLER_16_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13654_ clknet_leaf_42_clk _02283_ VGND VGND VPWR VPWR data_array.data1\[15\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10866_ net1022 net2894 net515 VGND VGND VPWR VPWR _02611_ sky130_fd_sc_hd__mux2_1
X_12605_ clknet_leaf_163_clk _01299_ VGND VGND VPWR VPWR tag_array.tag0\[0\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_13585_ clknet_leaf_111_clk _02214_ VGND VGND VPWR VPWR data_array.data0\[9\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_10797_ net1770 net1040 net502 VGND VGND VPWR VPWR _02542_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_171_3647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12536_ clknet_leaf_187_clk _01230_ VGND VGND VPWR VPWR tag_array.tag1\[11\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_173_904 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12467_ clknet_leaf_67_clk _01161_ VGND VGND VPWR VPWR data_array.data1\[9\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_14206_ clknet_leaf_221_clk _02835_ VGND VGND VPWR VPWR data_array.data0\[2\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_144_Right_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11418_ clknet_leaf_112_clk _00228_ VGND VGND VPWR VPWR data_array.data0\[0\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_12398_ clknet_leaf_222_clk _01092_ VGND VGND VPWR VPWR data_array.data0\[14\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_141_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14137_ clknet_leaf_53_clk _02766_ VGND VGND VPWR VPWR data_array.data0\[1\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
X_11349_ net898 net4578 net795 VGND VGND VPWR VPWR _03092_ sky130_fd_sc_hd__mux2_1
XFILLER_141_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14068_ clknet_leaf_84_clk _02697_ VGND VGND VPWR VPWR data_array.data1\[6\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_33_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05910_ data_array.rdata1\[26\] net828 net837 VGND VGND VPWR VPWR _03401_ sky130_fd_sc_hd__a21o_1
X_13019_ clknet_leaf_11_clk _01713_ VGND VGND VPWR VPWR data_array.data0\[3\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
X_06890_ _04180_ _04181_ VGND VGND VPWR VPWR _00004_ sky130_fd_sc_hd__or2_1
X_05841_ data_array.rdata1\[3\] net833 net842 VGND VGND VPWR VPWR _03355_ sky130_fd_sc_hd__a21o_1
XFILLER_94_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05772_ net3 fsm.tag_out1\[4\] VGND VGND VPWR VPWR _03289_ sky130_fd_sc_hd__and2b_1
X_08560_ net715 net4450 net585 VGND VGND VPWR VPWR _00328_ sky130_fd_sc_hd__mux2_1
XFILLER_47_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07511_ data_array.data1\[13\]\[6\] net1519 net1423 data_array.data1\[14\]\[6\] VGND
+ VGND VPWR VPWR _04746_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_18_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08491_ net824 _05550_ VGND VGND VPWR VPWR _05564_ sky130_fd_sc_hd__or2_1
XFILLER_81_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_5_1__f_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_5_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_07442_ data_array.data1\[12\]\[0\] net1366 net1272 data_array.data1\[15\]\[0\] _04682_
+ VGND VGND VPWR VPWR _04683_ sky130_fd_sc_hd__a221o_1
XFILLER_22_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07373_ net1217 _04615_ _04619_ net1169 VGND VGND VPWR VPWR _04621_ sky130_fd_sc_hd__a22o_1
XFILLER_22_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09112_ net1095 net2690 net574 VGND VGND VPWR VPWR _00866_ sky130_fd_sc_hd__mux2_1
XFILLER_13_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06324_ tag_array.tag0\[12\]\[12\] net1407 net1313 tag_array.tag0\[15\]\[12\] _03666_
+ VGND VGND VPWR VPWR _03667_ sky130_fd_sc_hd__a221o_1
XFILLER_30_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09043_ net807 _05574_ VGND VGND VPWR VPWR _05611_ sky130_fd_sc_hd__nand2_1
X_06255_ tag_array.tag0\[5\]\[6\] net1565 net1468 tag_array.tag0\[6\]\[6\] VGND VGND
+ VPWR VPWR _03604_ sky130_fd_sc_hd__a22o_1
XFILLER_108_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold410 data_array.data1\[0\]\[50\] VGND VGND VPWR VPWR net2061 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_111_Right_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06186_ _03540_ _03541_ VGND VGND VPWR VPWR _00182_ sky130_fd_sc_hd__or2_1
Xhold421 data_array.data1\[4\]\[6\] VGND VGND VPWR VPWR net2072 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold432 data_array.data1\[2\]\[45\] VGND VGND VPWR VPWR net2083 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold443 data_array.data1\[15\]\[17\] VGND VGND VPWR VPWR net2094 sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 data_array.data0\[2\]\[46\] VGND VGND VPWR VPWR net2105 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold465 data_array.data1\[4\]\[12\] VGND VGND VPWR VPWR net2116 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold476 data_array.data0\[6\]\[7\] VGND VGND VPWR VPWR net2127 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold487 data_array.data0\[4\]\[18\] VGND VGND VPWR VPWR net2138 sky130_fd_sc_hd__dlygate4sd3_1
Xhold498 data_array.data1\[0\]\[23\] VGND VGND VPWR VPWR net2149 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout901 _05524_ VGND VGND VPWR VPWR net901 sky130_fd_sc_hd__buf_1
X_09945_ net1048 net2126 net375 VGND VGND VPWR VPWR _01694_ sky130_fd_sc_hd__mux2_1
Xfanout912 _05518_ VGND VGND VPWR VPWR net912 sky130_fd_sc_hd__clkbuf_2
Xfanout923 _05514_ VGND VGND VPWR VPWR net923 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_70_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout934 _05508_ VGND VGND VPWR VPWR net934 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_70_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout945 net947 VGND VGND VPWR VPWR net945 sky130_fd_sc_hd__clkbuf_2
Xfanout956 net957 VGND VGND VPWR VPWR net956 sky130_fd_sc_hd__clkbuf_2
XFILLER_58_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout967 _05492_ VGND VGND VPWR VPWR net967 sky130_fd_sc_hd__dlymetal6s2s_1
X_09876_ net964 net3608 net384 VGND VGND VPWR VPWR _01626_ sky130_fd_sc_hd__mux2_1
XFILLER_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1110 data_array.data1\[3\]\[10\] VGND VGND VPWR VPWR net2761 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout978 net979 VGND VGND VPWR VPWR net978 sky130_fd_sc_hd__clkbuf_2
XFILLER_58_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout989 _05480_ VGND VGND VPWR VPWR net989 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1121 data_array.data1\[13\]\[51\] VGND VGND VPWR VPWR net2772 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_161_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1132 tag_array.tag0\[9\]\[14\] VGND VGND VPWR VPWR net2783 sky130_fd_sc_hd__dlygate4sd3_1
X_08827_ net1860 net938 net446 VGND VGND VPWR VPWR _00585_ sky130_fd_sc_hd__mux2_1
Xhold1143 data_array.data1\[9\]\[60\] VGND VGND VPWR VPWR net2794 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1154 tag_array.tag0\[13\]\[24\] VGND VGND VPWR VPWR net2805 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1165 data_array.data0\[5\]\[25\] VGND VGND VPWR VPWR net2816 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1176 data_array.data0\[10\]\[45\] VGND VGND VPWR VPWR net2827 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1187 data_array.data0\[1\]\[4\] VGND VGND VPWR VPWR net2838 sky130_fd_sc_hd__dlygate4sd3_1
X_08758_ net794 net3552 net451 VGND VGND VPWR VPWR _00517_ sky130_fd_sc_hd__mux2_1
Xhold1198 data_array.data1\[14\]\[63\] VGND VGND VPWR VPWR net2849 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07709_ data_array.data1\[9\]\[24\] net1585 net1489 data_array.data1\[10\]\[24\]
+ VGND VGND VPWR VPWR _04926_ sky130_fd_sc_hd__a22o_1
X_08689_ net1745 net766 net481 VGND VGND VPWR VPWR _00448_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_105_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10720_ net1094 net4367 net497 VGND VGND VPWR VPWR _02465_ sky130_fd_sc_hd__mux2_1
XFILLER_26_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1001 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10651_ net2140 net858 net469 VGND VGND VPWR VPWR _02396_ sky130_fd_sc_hd__mux2_1
XFILLER_55_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10582_ net879 net3543 net457 VGND VGND VPWR VPWR _02327_ sky130_fd_sc_hd__mux2_1
X_13370_ clknet_leaf_164_clk _02000_ VGND VGND VPWR VPWR tag_array.tag0\[2\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_142_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12321_ clknet_leaf_48_clk _00033_ VGND VGND VPWR VPWR data_array.rdata0\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_39_Left_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12252_ clknet_leaf_127_clk _01010_ VGND VGND VPWR VPWR tag_array.tag1\[14\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_163_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11203_ net963 net3199 net652 VGND VGND VPWR VPWR _02946_ sky130_fd_sc_hd__mux2_1
XFILLER_123_823 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12183_ clknet_leaf_162_clk _00991_ VGND VGND VPWR VPWR tag_array.tag0\[14\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_79_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11134_ net981 net4462 net541 VGND VGND VPWR VPWR _02877_ sky130_fd_sc_hd__mux2_1
XFILLER_122_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11065_ net2445 net1002 net331 VGND VGND VPWR VPWR _02808_ sky130_fd_sc_hd__mux2_1
XFILLER_122_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10016_ net1023 net3889 net556 VGND VGND VPWR VPWR _01765_ sky130_fd_sc_hd__mux2_1
XFILLER_77_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_48_Left_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11967_ clknet_leaf_244_clk _00775_ VGND VGND VPWR VPWR data_array.data0\[4\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13706_ clknet_leaf_253_clk _02335_ VGND VGND VPWR VPWR data_array.data1\[1\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_10918_ net1071 net4288 net535 VGND VGND VPWR VPWR _02663_ sky130_fd_sc_hd__mux2_1
XFILLER_60_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11898_ clknet_leaf_113_clk _00706_ VGND VGND VPWR VPWR data_array.data0\[5\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13637_ clknet_leaf_115_clk _02266_ VGND VGND VPWR VPWR data_array.data0\[9\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
X_10849_ net1090 net4364 net517 VGND VGND VPWR VPWR _02594_ sky130_fd_sc_hd__mux2_1
X_13568_ clknet_leaf_28_clk _02197_ VGND VGND VPWR VPWR tag_array.dirty1\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_57_Left_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12519_ clknet_leaf_233_clk _01213_ VGND VGND VPWR VPWR tag_array.tag1\[11\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13499_ clknet_leaf_29_clk _02128_ VGND VGND VPWR VPWR tag_array.dirty1\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_145_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06040_ fsm.tag_out0\[2\] net1120 _03483_ VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__a21o_1
XFILLER_154_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07991_ data_array.data1\[9\]\[50\] net1537 net1441 data_array.data1\[10\]\[50\]
+ VGND VGND VPWR VPWR _05182_ sky130_fd_sc_hd__a22o_1
XFILLER_140_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_7_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_7_0_clk sky130_fd_sc_hd__clkbuf_8
X_09730_ net766 net3939 net678 VGND VGND VPWR VPWR _01482_ sky130_fd_sc_hd__mux2_1
X_06942_ data_array.data0\[0\]\[18\] net1343 net1249 data_array.data0\[3\]\[18\] _04228_
+ VGND VGND VPWR VPWR _04229_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_66_Left_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09661_ net744 net2757 net612 VGND VGND VPWR VPWR _01413_ sky130_fd_sc_hd__mux2_1
X_06873_ data_array.data0\[13\]\[12\] net1579 net1483 data_array.data0\[14\]\[12\]
+ VGND VGND VPWR VPWR _04166_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_2_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08612_ net775 net3704 net516 VGND VGND VPWR VPWR _00371_ sky130_fd_sc_hd__mux2_1
X_05824_ _03237_ _03256_ _03339_ _03340_ VGND VGND VPWR VPWR _03341_ sky130_fd_sc_hd__or4_1
X_09592_ net983 net4595 net394 VGND VGND VPWR VPWR _01344_ sky130_fd_sc_hd__mux2_1
XFILLER_39_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08543_ net782 net2351 net581 VGND VGND VPWR VPWR _00311_ sky130_fd_sc_hd__mux2_1
X_05755_ fsm.tag_out1\[18\] net18 VGND VGND VPWR VPWR _03272_ sky130_fd_sc_hd__and2b_1
X_08474_ net1463 net1199 VGND VGND VPWR VPWR _05552_ sky130_fd_sc_hd__nand2_1
X_05686_ net13 fsm.tag_out0\[13\] VGND VGND VPWR VPWR _03203_ sky130_fd_sc_hd__xor2_1
XFILLER_168_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07425_ data_array.data0\[1\]\[62\] net1603 net1507 data_array.data0\[2\]\[62\] VGND
+ VGND VPWR VPWR _04668_ sky130_fd_sc_hd__a22o_1
XFILLER_126_1048 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_75_Left_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07356_ data_array.data0\[4\]\[56\] net1340 net1246 data_array.data0\[7\]\[56\] _04604_
+ VGND VGND VPWR VPWR _04605_ sky130_fd_sc_hd__a221o_1
XFILLER_164_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06307_ _03650_ _03651_ VGND VGND VPWR VPWR _00132_ sky130_fd_sc_hd__or2_1
X_07287_ data_array.data0\[9\]\[50\] net1540 net1444 data_array.data0\[10\]\[50\]
+ VGND VGND VPWR VPWR _04542_ sky130_fd_sc_hd__a22o_1
XFILLER_156_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06238_ tag_array.tag0\[0\]\[4\] net1371 net1277 tag_array.tag0\[3\]\[4\] _03588_
+ VGND VGND VPWR VPWR _03589_ sky130_fd_sc_hd__a221o_1
X_09026_ net2566 net921 net423 VGND VGND VPWR VPWR _00781_ sky130_fd_sc_hd__mux2_1
XFILLER_3_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold240 data_array.data1\[4\]\[15\] VGND VGND VPWR VPWR net1891 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_1043 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06169_ net29 net28 VGND VGND VPWR VPWR _03526_ sky130_fd_sc_hd__and2b_1
Xhold251 data_array.data1\[4\]\[4\] VGND VGND VPWR VPWR net1902 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 data_array.data0\[0\]\[61\] VGND VGND VPWR VPWR net1913 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold273 data_array.data0\[1\]\[46\] VGND VGND VPWR VPWR net1924 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold284 data_array.data0\[1\]\[21\] VGND VGND VPWR VPWR net1935 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 data_array.data1\[0\]\[41\] VGND VGND VPWR VPWR net1946 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout720 net721 VGND VGND VPWR VPWR net720 sky130_fd_sc_hd__clkbuf_2
Xfanout731 _05395_ VGND VGND VPWR VPWR net731 sky130_fd_sc_hd__buf_1
XFILLER_59_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09928_ net696 net4183 net604 VGND VGND VPWR VPWR _01678_ sky130_fd_sc_hd__mux2_1
Xfanout742 _05389_ VGND VGND VPWR VPWR net742 sky130_fd_sc_hd__clkbuf_2
Xfanout753 _05385_ VGND VGND VPWR VPWR net753 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout764 _05379_ VGND VGND VPWR VPWR net764 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_146_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout775 _05373_ VGND VGND VPWR VPWR net775 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout786 net788 VGND VGND VPWR VPWR net786 sky130_fd_sc_hd__clkbuf_2
X_09859_ net1033 net2067 net383 VGND VGND VPWR VPWR _01609_ sky130_fd_sc_hd__mux2_1
Xfanout797 net806 VGND VGND VPWR VPWR net797 sky130_fd_sc_hd__buf_4
XFILLER_86_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12870_ clknet_leaf_73_clk _01564_ VGND VGND VPWR VPWR data_array.data0\[12\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_142_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ clknet_leaf_175_clk _00629_ VGND VGND VPWR VPWR data_array.data0\[7\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11752_ clknet_leaf_47_clk _00560_ VGND VGND VPWR VPWR data_array.data0\[8\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_83_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ net2235 net906 net478 VGND VGND VPWR VPWR _02448_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_120_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14471_ clknet_leaf_17_clk _03094_ VGND VGND VPWR VPWR data_array.data1\[7\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11683_ clknet_leaf_189_clk _00491_ VGND VGND VPWR VPWR tag_array.tag1\[1\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_13422_ clknet_leaf_88_clk _02052_ VGND VGND VPWR VPWR data_array.data1\[8\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
X_10634_ net2281 net924 net466 VGND VGND VPWR VPWR _02379_ sky130_fd_sc_hd__mux2_1
XFILLER_155_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13353_ clknet_leaf_115_clk _01983_ VGND VGND VPWR VPWR data_array.data0\[10\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
X_10565_ net944 net3898 net453 VGND VGND VPWR VPWR _02310_ sky130_fd_sc_hd__mux2_1
XFILLER_127_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12304_ clknet_leaf_97_clk _01062_ VGND VGND VPWR VPWR tag_array.tag1\[12\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_13284_ clknet_leaf_237_clk _01914_ VGND VGND VPWR VPWR data_array.data0\[11\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
X_10496_ net962 net3569 net346 VGND VGND VPWR VPWR _02241_ sky130_fd_sc_hd__mux2_1
XFILLER_170_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12235_ clknet_leaf_147_clk _00164_ VGND VGND VPWR VPWR fsm.tag_out1\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_151_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_166_3546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12166_ clknet_leaf_159_clk _00974_ VGND VGND VPWR VPWR tag_array.tag0\[13\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_11117_ net1050 net4217 net549 VGND VGND VPWR VPWR _02860_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_183_3871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_3882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12097_ clknet_leaf_43_clk _00905_ VGND VGND VPWR VPWR data_array.data1\[14\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_127_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11048_ net1773 net1068 net335 VGND VGND VPWR VPWR _02791_ sky130_fd_sc_hd__mux2_1
XFILLER_76_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput8 cpu_addr[16] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_2
XFILLER_52_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12999_ clknet_leaf_50_clk _01693_ VGND VGND VPWR VPWR data_array.data0\[3\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07210_ data_array.data0\[9\]\[43\] net1569 net1473 data_array.data0\[10\]\[43\]
+ VGND VGND VPWR VPWR _04472_ sky130_fd_sc_hd__a22o_1
X_08190_ net1644 _03347_ _05358_ _05357_ VGND VGND VPWR VPWR _05360_ sky130_fd_sc_hd__a31o_1
X_07141_ net1635 _04403_ _04407_ net1209 VGND VGND VPWR VPWR _04410_ sky130_fd_sc_hd__a22o_1
XFILLER_146_723 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07072_ data_array.data0\[12\]\[30\] net1391 net1297 data_array.data0\[15\]\[30\]
+ _04346_ VGND VGND VPWR VPWR _04347_ sky130_fd_sc_hd__a221o_1
Xoutput301 net301 VGND VGND VPWR VPWR mem_wdata[44] sky130_fd_sc_hd__buf_2
XFILLER_105_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput312 net312 VGND VGND VPWR VPWR mem_wdata[54] sky130_fd_sc_hd__buf_2
X_06023_ net1164 net1 VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__and2_1
Xoutput323 net323 VGND VGND VPWR VPWR mem_wdata[6] sky130_fd_sc_hd__buf_2
XFILLER_99_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07974_ data_array.data1\[12\]\[48\] net1393 net1299 data_array.data1\[15\]\[48\]
+ _05166_ VGND VGND VPWR VPWR _05167_ sky130_fd_sc_hd__a221o_1
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09713_ net736 net2926 net609 VGND VGND VPWR VPWR _01465_ sky130_fd_sc_hd__mux2_1
X_06925_ data_array.data0\[12\]\[17\] net1338 net1244 data_array.data0\[15\]\[17\]
+ _04212_ VGND VGND VPWR VPWR _04213_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_87_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09644_ net712 net4008 net615 VGND VGND VPWR VPWR _01396_ sky130_fd_sc_hd__mux2_1
X_06856_ net1183 _04145_ _04149_ net1231 VGND VGND VPWR VPWR _04151_ sky130_fd_sc_hd__a22o_1
XFILLER_55_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05807_ _03174_ _03175_ _03322_ _03323_ VGND VGND VPWR VPWR _03324_ sky130_fd_sc_hd__or4_1
X_09575_ net1048 net3534 net399 VGND VGND VPWR VPWR _01327_ sky130_fd_sc_hd__mux2_1
XFILLER_71_927 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06787_ data_array.data0\[1\]\[4\] net1581 net1485 data_array.data0\[2\]\[4\] VGND
+ VGND VPWR VPWR _04088_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_65_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08526_ net821 net812 net854 _05587_ VGND VGND VPWR VPWR _05589_ sky130_fd_sc_hd__or4b_1
XFILLER_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05738_ _03245_ _03246_ _03254_ _03244_ VGND VGND VPWR VPWR _03255_ sky130_fd_sc_hd__or4b_1
X_08457_ net156 net91 net1645 VGND VGND VPWR VPWR _05541_ sky130_fd_sc_hd__mux2_1
XFILLER_23_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05669_ _03182_ _03183_ _03184_ _03185_ VGND VGND VPWR VPWR _03186_ sky130_fd_sc_hd__or4_1
X_07408_ data_array.data0\[13\]\[61\] net1553 net1457 data_array.data0\[14\]\[61\]
+ VGND VGND VPWR VPWR _04652_ sky130_fd_sc_hd__a22o_1
X_08388_ net130 net65 net1641 VGND VGND VPWR VPWR _05495_ sky130_fd_sc_hd__mux2_1
XFILLER_149_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07339_ net1621 _04583_ _04587_ net1195 VGND VGND VPWR VPWR _04590_ sky130_fd_sc_hd__a22o_1
XFILLER_167_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10350_ net699 net3642 net592 VGND VGND VPWR VPWR _02097_ sky130_fd_sc_hd__mux2_1
XFILLER_152_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09009_ net2129 net988 net422 VGND VGND VPWR VPWR _00764_ sky130_fd_sc_hd__mux2_1
XFILLER_152_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10281_ net2921 net1039 net635 VGND VGND VPWR VPWR _02028_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_148_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_758 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12020_ clknet_leaf_71_clk _00828_ VGND VGND VPWR VPWR data_array.data0\[6\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1504 net1517 VGND VGND VPWR VPWR net1504 sky130_fd_sc_hd__clkbuf_2
Xfanout1515 net1516 VGND VGND VPWR VPWR net1515 sky130_fd_sc_hd__buf_2
Xfanout1526 net1530 VGND VGND VPWR VPWR net1526 sky130_fd_sc_hd__clkbuf_4
Xfanout1537 net1539 VGND VGND VPWR VPWR net1537 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_144_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout550 net553 VGND VGND VPWR VPWR net550 sky130_fd_sc_hd__clkbuf_4
Xfanout1548 net1549 VGND VGND VPWR VPWR net1548 sky130_fd_sc_hd__clkbuf_4
Xfanout1559 net1560 VGND VGND VPWR VPWR net1559 sky130_fd_sc_hd__clkbuf_4
Xfanout561 net563 VGND VGND VPWR VPWR net561 sky130_fd_sc_hd__clkbuf_8
Xfanout572 _05592_ VGND VGND VPWR VPWR net572 sky130_fd_sc_hd__clkbuf_4
XFILLER_19_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout583 net584 VGND VGND VPWR VPWR net583 sky130_fd_sc_hd__buf_2
X_13971_ clknet_leaf_35_clk _02600_ VGND VGND VPWR VPWR data_array.data1\[5\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_161_3454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout594 _05589_ VGND VGND VPWR VPWR net594 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_161_3465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12922_ clknet_leaf_245_clk _01616_ VGND VGND VPWR VPWR data_array.data0\[13\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_46_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_122_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12853_ clknet_leaf_226_clk _01547_ VGND VGND VPWR VPWR data_array.data0\[12\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_92_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11804_ clknet_leaf_270_clk _00612_ VGND VGND VPWR VPWR data_array.data0\[7\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12784_ clknet_leaf_32_clk _01478_ VGND VGND VPWR VPWR tag_array.tag1\[10\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_11735_ clknet_leaf_261_clk _00543_ VGND VGND VPWR VPWR data_array.data0\[8\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14454_ clknet_leaf_74_clk _03077_ VGND VGND VPWR VPWR data_array.data1\[7\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_159_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11666_ clknet_leaf_132_clk _00474_ VGND VGND VPWR VPWR tag_array.tag1\[1\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13405_ clknet_leaf_263_clk _02035_ VGND VGND VPWR VPWR data_array.data1\[8\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_10617_ net3928 net995 net471 VGND VGND VPWR VPWR _02362_ sky130_fd_sc_hd__mux2_1
X_14385_ clknet_leaf_258_clk _03008_ VGND VGND VPWR VPWR data_array.data1\[10\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
X_11597_ clknet_leaf_133_clk _00405_ VGND VGND VPWR VPWR tag_array.tag1\[4\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_13336_ clknet_leaf_22_clk _01966_ VGND VGND VPWR VPWR data_array.data0\[10\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
X_10548_ net1014 net3887 net462 VGND VGND VPWR VPWR _02293_ sky130_fd_sc_hd__mux2_1
XFILLER_182_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13267_ clknet_leaf_124_clk _01897_ VGND VGND VPWR VPWR data_array.data0\[11\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
X_10479_ net1029 net3197 net350 VGND VGND VPWR VPWR _02224_ sky130_fd_sc_hd__mux2_1
XFILLER_68_1071 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12218_ clknet_5_29__leaf_clk _00156_ VGND VGND VPWR VPWR fsm.tag_out1\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_170_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13198_ clknet_leaf_256_clk _00092_ VGND VGND VPWR VPWR data_array.rdata1\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_151_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_1074 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12149_ clknet_leaf_153_clk _00957_ VGND VGND VPWR VPWR tag_array.tag0\[13\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_69_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1709 tag_array.tag0\[2\]\[22\] VGND VGND VPWR VPWR net3360 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06710_ tag_array.tag1\[5\]\[22\] net1552 net1456 tag_array.tag1\[6\]\[22\] VGND
+ VGND VPWR VPWR _04018_ sky130_fd_sc_hd__a22o_1
XFILLER_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07690_ data_array.data1\[4\]\[22\] net1341 net1247 data_array.data1\[7\]\[22\] _04908_
+ VGND VGND VPWR VPWR _04909_ sky130_fd_sc_hd__a221o_1
XFILLER_37_467 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06641_ tag_array.tag1\[0\]\[16\] net1417 net1323 tag_array.tag1\[3\]\[16\] _03954_
+ VGND VGND VPWR VPWR _03955_ sky130_fd_sc_hd__a221o_1
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09360_ net961 net2307 net404 VGND VGND VPWR VPWR _01113_ sky130_fd_sc_hd__mux2_1
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06572_ tag_array.tag1\[13\]\[10\] net1595 net1499 tag_array.tag1\[14\]\[10\] VGND
+ VGND VPWR VPWR _03892_ sky130_fd_sc_hd__a22o_1
X_08311_ net1129 _05443_ VGND VGND VPWR VPWR _05444_ sky130_fd_sc_hd__and2_1
XFILLER_177_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09291_ net714 net3378 net561 VGND VGND VPWR VPWR _01045_ sky130_fd_sc_hd__mux2_1
XFILLER_36_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_13 _03132_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_846 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08242_ net1650 net1163 net16 VGND VGND VPWR VPWR _05396_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_60_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_24 _05367_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_35 net385 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_46 net594 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_57 net1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08173_ lru_array.lru_mem\[1\] net1563 net1467 lru_array.lru_mem\[2\] VGND VGND VPWR
+ VPWR _05348_ sky130_fd_sc_hd__a22o_1
XANTENNA_68 net1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_79 net417 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07124_ data_array.data0\[5\]\[35\] net1537 net1441 data_array.data0\[6\]\[35\] VGND
+ VGND VPWR VPWR _04394_ sky130_fd_sc_hd__a22o_1
XFILLER_137_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07055_ _04330_ _04331_ VGND VGND VPWR VPWR _00020_ sky130_fd_sc_hd__or2_2
X_06006_ data_array.rdata1\[58\] net830 net840 VGND VGND VPWR VPWR _03465_ sky130_fd_sc_hd__a21o_1
XFILLER_115_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput175 net175 VGND VGND VPWR VPWR cpu_rdata[19] sky130_fd_sc_hd__buf_6
XFILLER_82_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput186 net186 VGND VGND VPWR VPWR cpu_rdata[29] sky130_fd_sc_hd__clkbuf_4
Xhold2900 tag_array.tag1\[12\]\[9\] VGND VGND VPWR VPWR net4551 sky130_fd_sc_hd__dlygate4sd3_1
Xoutput197 net197 VGND VGND VPWR VPWR cpu_rdata[39] sky130_fd_sc_hd__clkbuf_4
XFILLER_88_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2911 data_array.data0\[7\]\[50\] VGND VGND VPWR VPWR net4562 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2922 data_array.data0\[12\]\[23\] VGND VGND VPWR VPWR net4573 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_87_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2933 tag_array.tag0\[4\]\[6\] VGND VGND VPWR VPWR net4584 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2944 data_array.data0\[15\]\[32\] VGND VGND VPWR VPWR net4595 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2955 data_array.data0\[10\]\[55\] VGND VGND VPWR VPWR net4606 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2966 data_array.data1\[3\]\[25\] VGND VGND VPWR VPWR net4617 sky130_fd_sc_hd__dlygate4sd3_1
X_07957_ _05150_ _05151_ VGND VGND VPWR VPWR _00104_ sky130_fd_sc_hd__or2_1
X_06908_ data_array.data0\[1\]\[15\] net1582 net1486 data_array.data0\[2\]\[15\] VGND
+ VGND VPWR VPWR _04198_ sky130_fd_sc_hd__a22o_1
X_07888_ data_array.data1\[0\]\[40\] net1415 net1321 data_array.data1\[3\]\[40\] _05088_
+ VGND VGND VPWR VPWR _05089_ sky130_fd_sc_hd__a221o_1
XFILLER_55_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09627_ net781 net3117 net615 VGND VGND VPWR VPWR _01379_ sky130_fd_sc_hd__mux2_1
X_06839_ data_array.data0\[4\]\[9\] net1389 net1295 data_array.data0\[7\]\[9\] _04134_
+ VGND VGND VPWR VPWR _04135_ sky130_fd_sc_hd__a221o_1
X_09558_ net694 net2607 net620 VGND VGND VPWR VPWR _01311_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08509_ net1703 net611 VGND VGND VPWR VPWR _00298_ sky130_fd_sc_hd__nand2b_1
XFILLER_12_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09489_ net771 net4157 net626 VGND VGND VPWR VPWR _01242_ sky130_fd_sc_hd__mux2_1
XFILLER_11_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11520_ clknet_leaf_103_clk _00328_ VGND VGND VPWR VPWR tag_array.tag1\[9\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11451_ clknet_leaf_125_clk _00261_ VGND VGND VPWR VPWR data_array.data0\[0\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10402_ net2257 net1044 net664 VGND VGND VPWR VPWR _02148_ sky130_fd_sc_hd__mux2_1
XFILLER_183_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14170_ clknet_leaf_15_clk _02799_ VGND VGND VPWR VPWR data_array.data0\[2\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_11382_ net164 VGND VGND VPWR VPWR _00192_ sky130_fd_sc_hd__inv_2
XFILLER_165_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_12_Left_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13121_ clknet_leaf_144_clk _01815_ VGND VGND VPWR VPWR tag_array.tag0\[3\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_10333_ net768 net4590 net591 VGND VGND VPWR VPWR _02080_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_115_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13052_ clknet_leaf_36_clk _01746_ VGND VGND VPWR VPWR data_array.data1\[13\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_106_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10264_ net2130 net1107 net633 VGND VGND VPWR VPWR _02011_ sky130_fd_sc_hd__mux2_1
XFILLER_97_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12003_ clknet_leaf_224_clk _00811_ VGND VGND VPWR VPWR data_array.data0\[6\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1301 net1305 VGND VGND VPWR VPWR net1301 sky130_fd_sc_hd__clkbuf_4
X_10195_ net1026 net3858 net357 VGND VGND VPWR VPWR _01942_ sky130_fd_sc_hd__mux2_1
Xfanout1312 net1328 VGND VGND VPWR VPWR net1312 sky130_fd_sc_hd__buf_2
Xfanout1323 net1327 VGND VGND VPWR VPWR net1323 sky130_fd_sc_hd__clkbuf_4
Xfanout1334 net1376 VGND VGND VPWR VPWR net1334 sky130_fd_sc_hd__buf_2
XFILLER_87_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1345 net1352 VGND VGND VPWR VPWR net1345 sky130_fd_sc_hd__clkbuf_4
XFILLER_38_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1356 net1358 VGND VGND VPWR VPWR net1356 sky130_fd_sc_hd__clkbuf_4
Xfanout1367 net1370 VGND VGND VPWR VPWR net1367 sky130_fd_sc_hd__clkbuf_2
XFILLER_4_1013 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout380 net381 VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__buf_4
Xfanout1378 net1383 VGND VGND VPWR VPWR net1378 sky130_fd_sc_hd__clkbuf_4
Xfanout391 net392 VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__buf_4
Xfanout1389 net1392 VGND VGND VPWR VPWR net1389 sky130_fd_sc_hd__clkbuf_4
XFILLER_93_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13954_ clknet_leaf_201_clk _02583_ VGND VGND VPWR VPWR data_array.data1\[4\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
X_12905_ clknet_leaf_60_clk _01599_ VGND VGND VPWR VPWR data_array.data0\[13\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_938 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_194_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_194_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13885_ clknet_leaf_5_clk _02514_ VGND VGND VPWR VPWR data_array.data1\[3\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_98_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12836_ clknet_leaf_71_clk _01530_ VGND VGND VPWR VPWR data_array.data0\[12\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_178_3781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12767_ clknet_leaf_105_clk _01461_ VGND VGND VPWR VPWR tag_array.tag0\[6\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11718_ clknet_leaf_158_clk _00526_ VGND VGND VPWR VPWR tag_array.tag0\[9\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_12698_ clknet_leaf_157_clk _01392_ VGND VGND VPWR VPWR tag_array.tag0\[8\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_159_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14437_ clknet_leaf_229_clk _03060_ VGND VGND VPWR VPWR data_array.data1\[7\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput11 cpu_addr[19] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dlymetal6s2s_1
X_11649_ clknet_leaf_98_clk _00457_ VGND VGND VPWR VPWR tag_array.tag1\[2\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput22 cpu_addr[29] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_2
XFILLER_156_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput33 cpu_read VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_1
Xinput44 cpu_wdata[19] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_1
X_14368_ clknet_leaf_19_clk _02991_ VGND VGND VPWR VPWR data_array.data1\[10\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput55 cpu_wdata[29] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_1
XFILLER_183_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput66 cpu_wdata[39] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_1
Xhold806 data_array.data0\[0\]\[32\] VGND VGND VPWR VPWR net2457 sky130_fd_sc_hd__dlygate4sd3_1
Xinput77 cpu_wdata[49] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_1
Xhold817 data_array.data0\[1\]\[39\] VGND VGND VPWR VPWR net2468 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_183_692 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold828 tag_array.tag1\[11\]\[5\] VGND VGND VPWR VPWR net2479 sky130_fd_sc_hd__dlygate4sd3_1
X_13319_ clknet_leaf_30_clk _01949_ VGND VGND VPWR VPWR data_array.data0\[10\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput88 cpu_wdata[59] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__clkbuf_1
Xhold839 data_array.data0\[15\]\[35\] VGND VGND VPWR VPWR net2490 sky130_fd_sc_hd__dlygate4sd3_1
Xinput99 mem_rdata[0] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_1
X_14299_ clknet_leaf_67_clk _02928_ VGND VGND VPWR VPWR data_array.data1\[11\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_171_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2207 data_array.data0\[10\]\[21\] VGND VGND VPWR VPWR net3858 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08860_ net1064 net4256 net439 VGND VGND VPWR VPWR _00617_ sky130_fd_sc_hd__mux2_1
Xhold2218 data_array.data1\[15\]\[33\] VGND VGND VPWR VPWR net3869 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2229 tag_array.tag0\[12\]\[5\] VGND VGND VPWR VPWR net3880 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_36_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1506 data_array.data1\[10\]\[40\] VGND VGND VPWR VPWR net3157 sky130_fd_sc_hd__dlygate4sd3_1
X_07811_ data_array.data1\[4\]\[33\] net1397 net1303 data_array.data1\[7\]\[33\] _05018_
+ VGND VGND VPWR VPWR _05019_ sky130_fd_sc_hd__a221o_1
Xhold1517 data_array.data1\[7\]\[61\] VGND VGND VPWR VPWR net3168 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08791_ net1778 net1081 net448 VGND VGND VPWR VPWR _00549_ sky130_fd_sc_hd__mux2_1
XFILLER_85_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1528 data_array.data0\[5\]\[62\] VGND VGND VPWR VPWR net3179 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1539 data_array.data1\[10\]\[45\] VGND VGND VPWR VPWR net3190 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07742_ data_array.data1\[13\]\[27\] net1549 net1453 data_array.data1\[14\]\[27\]
+ VGND VGND VPWR VPWR _04956_ sky130_fd_sc_hd__a22o_1
XFILLER_42_1074 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07673_ data_array.data1\[8\]\[21\] net1365 net1271 data_array.data1\[11\]\[21\]
+ _04892_ VGND VGND VPWR VPWR _04893_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_185_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_185_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_93_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09412_ net1017 net4109 net582 VGND VGND VPWR VPWR _01165_ sky130_fd_sc_hd__mux2_1
X_06624_ net1625 _03933_ _03937_ net1199 VGND VGND VPWR VPWR _03940_ sky130_fd_sc_hd__a22o_1
XFILLER_179_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09343_ net1028 net4284 net408 VGND VGND VPWR VPWR _01096_ sky130_fd_sc_hd__mux2_1
XFILLER_12_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06555_ tag_array.tag1\[12\]\[8\] net1417 net1323 tag_array.tag1\[15\]\[8\] _03876_
+ VGND VGND VPWR VPWR _03877_ sky130_fd_sc_hd__a221o_1
XFILLER_179_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_158_Right_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09274_ net783 net3633 net557 VGND VGND VPWR VPWR _01028_ sky130_fd_sc_hd__mux2_1
X_06486_ tag_array.tag1\[5\]\[2\] net1541 net1445 tag_array.tag1\[6\]\[2\] VGND VGND
+ VPWR VPWR _03814_ sky130_fd_sc_hd__a22o_1
XFILLER_178_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08225_ fsm.tag_out1\[10\] net817 net809 fsm.tag_out0\[10\] _05384_ VGND VGND VPWR
+ VPWR _05385_ sky130_fd_sc_hd__a221o_1
XFILLER_21_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08156_ tag_array.dirty0\[13\] net1594 net1498 tag_array.dirty0\[14\] VGND VGND VPWR
+ VPWR _05332_ sky130_fd_sc_hd__a22o_1
XFILLER_162_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07107_ data_array.data0\[4\]\[33\] net1396 net1302 data_array.data0\[7\]\[33\] _04378_
+ VGND VGND VPWR VPWR _04379_ sky130_fd_sc_hd__a221o_1
XFILLER_180_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08087_ net1622 _05263_ _05267_ net1196 VGND VGND VPWR VPWR _05270_ sky130_fd_sc_hd__a22o_1
XFILLER_164_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07038_ data_array.data0\[13\]\[27\] net1538 net1442 data_array.data0\[14\]\[27\]
+ VGND VGND VPWR VPWR _04316_ sky130_fd_sc_hd__a22o_1
XFILLER_103_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2730 tag_array.dirty1\[6\] VGND VGND VPWR VPWR net4381 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_110_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2741 tag_array.tag0\[15\]\[4\] VGND VGND VPWR VPWR net4392 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2752 data_array.data1\[7\]\[54\] VGND VGND VPWR VPWR net4403 sky130_fd_sc_hd__dlygate4sd3_1
X_08989_ net2174 net1069 net424 VGND VGND VPWR VPWR _00744_ sky130_fd_sc_hd__mux2_1
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2763 data_array.data0\[14\]\[43\] VGND VGND VPWR VPWR net4414 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2774 tag_array.tag1\[5\]\[15\] VGND VGND VPWR VPWR net4425 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2785 tag_array.tag0\[13\]\[10\] VGND VGND VPWR VPWR net4436 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2796 data_array.data0\[7\]\[28\] VGND VGND VPWR VPWR net4447 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10951_ net937 net4412 net531 VGND VGND VPWR VPWR _02696_ sky130_fd_sc_hd__mux2_1
XFILLER_29_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_176_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_176_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_44_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13670_ clknet_leaf_67_clk _02299_ VGND VGND VPWR VPWR data_array.data1\[15\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_44_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10882_ net958 net4166 net521 VGND VGND VPWR VPWR _02627_ sky130_fd_sc_hd__mux2_1
XFILLER_43_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12621_ clknet_leaf_46_clk _01315_ VGND VGND VPWR VPWR data_array.data0\[15\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_139_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_125_Right_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_156_3353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12552_ clknet_leaf_158_clk _01246_ VGND VGND VPWR VPWR tag_array.tag0\[11\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_129_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11503_ clknet_leaf_32_clk _00311_ VGND VGND VPWR VPWR tag_array.tag1\[9\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_184_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12483_ clknet_leaf_259_clk _01177_ VGND VGND VPWR VPWR data_array.data1\[9\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_20_Left_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14222_ clknet_leaf_268_clk _02851_ VGND VGND VPWR VPWR data_array.data1\[12\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_11434_ clknet_leaf_175_clk _00244_ VGND VGND VPWR VPWR data_array.data0\[0\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_134_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14153_ clknet_leaf_262_clk _02782_ VGND VGND VPWR VPWR data_array.data0\[2\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_100_clk clknet_5_24__leaf_clk VGND VGND VPWR VPWR clknet_leaf_100_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11365_ net1646 net4159 net603 VGND VGND VPWR VPWR _03108_ sky130_fd_sc_hd__mux2_1
XFILLER_138_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13104_ clknet_leaf_21_clk _01798_ VGND VGND VPWR VPWR data_array.data1\[13\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_180_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10316_ net2041 net899 net633 VGND VGND VPWR VPWR _02063_ sky130_fd_sc_hd__mux2_1
X_14084_ clknet_leaf_120_clk _02713_ VGND VGND VPWR VPWR data_array.data1\[6\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11296_ net1110 net3824 net799 VGND VGND VPWR VPWR _03039_ sky130_fd_sc_hd__mux2_1
XFILLER_140_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13035_ clknet_leaf_241_clk _01729_ VGND VGND VPWR VPWR data_array.data0\[3\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
X_10247_ net754 net3430 net597 VGND VGND VPWR VPWR _01994_ sky130_fd_sc_hd__mux2_1
XFILLER_65_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1120 _03478_ VGND VGND VPWR VPWR net1120 sky130_fd_sc_hd__clkbuf_4
Xfanout1131 net1133 VGND VGND VPWR VPWR net1131 sky130_fd_sc_hd__buf_2
Xfanout1142 net1143 VGND VGND VPWR VPWR net1142 sky130_fd_sc_hd__buf_4
XFILLER_120_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10178_ net1092 net3854 net359 VGND VGND VPWR VPWR _01925_ sky130_fd_sc_hd__mux2_1
XFILLER_67_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1153 net1154 VGND VGND VPWR VPWR net1153 sky130_fd_sc_hd__clkbuf_4
Xfanout1164 net262 VGND VGND VPWR VPWR net1164 sky130_fd_sc_hd__clkbuf_2
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1175 _03526_ VGND VGND VPWR VPWR net1175 sky130_fd_sc_hd__clkbuf_4
Xfanout1186 net1187 VGND VGND VPWR VPWR net1186 sky130_fd_sc_hd__clkbuf_4
Xfanout1197 net1198 VGND VGND VPWR VPWR net1197 sky130_fd_sc_hd__clkbuf_2
XFILLER_47_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13937_ clknet_leaf_258_clk _02566_ VGND VGND VPWR VPWR data_array.data1\[4\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_167_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_167_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13868_ clknet_leaf_116_clk _02497_ VGND VGND VPWR VPWR data_array.data1\[3\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
X_12819_ clknet_leaf_167_clk _01513_ VGND VGND VPWR VPWR tag_array.tag1\[0\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_13799_ clknet_leaf_41_clk _02428_ VGND VGND VPWR VPWR data_array.data1\[2\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_06340_ _03680_ _03681_ VGND VGND VPWR VPWR _00135_ sky130_fd_sc_hd__or2_1
XFILLER_31_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06271_ tag_array.tag0\[4\]\[7\] net1418 net1324 tag_array.tag0\[7\]\[7\] _03618_
+ VGND VGND VPWR VPWR _03619_ sky130_fd_sc_hd__a221o_1
XFILLER_176_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08010_ net1189 _05193_ _05197_ net1615 VGND VGND VPWR VPWR _05200_ sky130_fd_sc_hd__a22o_1
XFILLER_147_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold603 data_array.data0\[0\]\[43\] VGND VGND VPWR VPWR net2254 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold614 data_array.data0\[2\]\[61\] VGND VGND VPWR VPWR net2265 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold625 data_array.data0\[1\]\[42\] VGND VGND VPWR VPWR net2276 sky130_fd_sc_hd__dlygate4sd3_1
Xhold636 data_array.data1\[2\]\[38\] VGND VGND VPWR VPWR net2287 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold647 data_array.data1\[0\]\[46\] VGND VGND VPWR VPWR net2298 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_94_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold658 data_array.data1\[9\]\[17\] VGND VGND VPWR VPWR net2309 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09961_ net986 net3166 net376 VGND VGND VPWR VPWR _01710_ sky130_fd_sc_hd__mux2_1
Xhold669 data_array.data0\[0\]\[10\] VGND VGND VPWR VPWR net2320 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08912_ net856 net4139 net437 VGND VGND VPWR VPWR _00669_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09892_ net902 net4066 net381 VGND VGND VPWR VPWR _01642_ sky130_fd_sc_hd__mux2_1
Xhold2004 tag_array.tag0\[3\]\[2\] VGND VGND VPWR VPWR net3655 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2015 data_array.data1\[7\]\[12\] VGND VGND VPWR VPWR net3666 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2026 data_array.data1\[14\]\[55\] VGND VGND VPWR VPWR net3677 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2037 data_array.data0\[7\]\[36\] VGND VGND VPWR VPWR net3688 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08843_ net2327 net872 net446 VGND VGND VPWR VPWR _00601_ sky130_fd_sc_hd__mux2_1
Xhold1303 data_array.data0\[12\]\[40\] VGND VGND VPWR VPWR net2954 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2048 data_array.data1\[10\]\[54\] VGND VGND VPWR VPWR net3699 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2059 data_array.data1\[3\]\[32\] VGND VGND VPWR VPWR net3710 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1314 data_array.data0\[12\]\[3\] VGND VGND VPWR VPWR net2965 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1325 tag_array.tag0\[12\]\[6\] VGND VGND VPWR VPWR net2976 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1336 data_array.data1\[13\]\[10\] VGND VGND VPWR VPWR net2987 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1347 data_array.data1\[11\]\[58\] VGND VGND VPWR VPWR net2998 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08774_ net726 net4476 net452 VGND VGND VPWR VPWR _00533_ sky130_fd_sc_hd__mux2_1
X_05986_ net145 net1150 _03450_ _03451_ VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__a22o_1
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1358 data_array.data0\[9\]\[13\] VGND VGND VPWR VPWR net3009 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1369 data_array.data0\[15\]\[8\] VGND VGND VPWR VPWR net3020 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07725_ net1213 _04935_ _04939_ net1165 VGND VGND VPWR VPWR _04941_ sky130_fd_sc_hd__a22o_1
XFILLER_84_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_158_clk clknet_5_28__leaf_clk VGND VGND VPWR VPWR clknet_leaf_158_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07656_ data_array.data1\[1\]\[19\] net1584 net1488 data_array.data1\[2\]\[19\] VGND
+ VGND VPWR VPWR _04878_ sky130_fd_sc_hd__a22o_1
XFILLER_53_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06607_ tag_array.tag1\[5\]\[13\] net1611 net1515 tag_array.tag1\[6\]\[13\] VGND
+ VGND VPWR VPWR _03924_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07587_ data_array.data1\[0\]\[13\] net1360 net1266 data_array.data1\[3\]\[13\] _04814_
+ VGND VGND VPWR VPWR _04815_ sky130_fd_sc_hd__a221o_1
XFILLER_40_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09326_ net1097 net4320 net406 VGND VGND VPWR VPWR _01079_ sky130_fd_sc_hd__mux2_1
X_06538_ _03860_ _03861_ VGND VGND VPWR VPWR _00177_ sky130_fd_sc_hd__or2_1
XFILLER_21_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09257_ net751 net3267 net577 VGND VGND VPWR VPWR _01011_ sky130_fd_sc_hd__mux2_1
X_06469_ tag_array.tag1\[4\]\[0\] net1385 net1291 tag_array.tag1\[7\]\[0\] _03798_
+ VGND VGND VPWR VPWR _03799_ sky130_fd_sc_hd__a221o_1
XFILLER_182_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08208_ net774 net2329 net798 VGND VGND VPWR VPWR _00200_ sky130_fd_sc_hd__mux2_1
XFILLER_126_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_151_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09188_ net727 net2614 net628 VGND VGND VPWR VPWR _00942_ sky130_fd_sc_hd__mux2_1
XFILLER_182_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08139_ data_array.data1\[8\]\[63\] net1363 net1269 data_array.data1\[11\]\[63\]
+ _05316_ VGND VGND VPWR VPWR _05317_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_75_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11150_ net919 net3299 net549 VGND VGND VPWR VPWR _02893_ sky130_fd_sc_hd__mux2_1
XFILLER_49_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1069 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10101_ net2179 net718 net638 VGND VGND VPWR VPWR _01850_ sky130_fd_sc_hd__mux2_1
XFILLER_108_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11081_ net3051 net936 net334 VGND VGND VPWR VPWR _02824_ sky130_fd_sc_hd__mux2_1
XFILLER_68_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10032_ net959 net4345 net562 VGND VGND VPWR VPWR _01781_ sky130_fd_sc_hd__mux2_1
XFILLER_102_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2560 tag_array.tag1\[7\]\[1\] VGND VGND VPWR VPWR net4211 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2571 data_array.data0\[9\]\[32\] VGND VGND VPWR VPWR net4222 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2582 data_array.data0\[11\]\[57\] VGND VGND VPWR VPWR net4233 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2593 data_array.data0\[3\]\[33\] VGND VGND VPWR VPWR net4244 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_63_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1870 tag_array.tag0\[10\]\[17\] VGND VGND VPWR VPWR net3521 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1881 data_array.data0\[13\]\[40\] VGND VGND VPWR VPWR net3532 sky130_fd_sc_hd__dlygate4sd3_1
X_11983_ clknet_leaf_236_clk _00791_ VGND VGND VPWR VPWR data_array.data0\[4\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1892 data_array.data1\[15\]\[58\] VGND VGND VPWR VPWR net3543 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_16_223 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13722_ clknet_leaf_18_clk _02351_ VGND VGND VPWR VPWR data_array.data1\[1\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_158_3404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10934_ net1004 net2908 net527 VGND VGND VPWR VPWR _02679_ sky130_fd_sc_hd__mux2_1
XFILLER_140_50 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13653_ clknet_leaf_199_clk _02282_ VGND VGND VPWR VPWR data_array.data1\[15\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_44_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10865_ net1024 net4438 net517 VGND VGND VPWR VPWR _02610_ sky130_fd_sc_hd__mux2_1
XFILLER_31_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12604_ clknet_leaf_165_clk _01298_ VGND VGND VPWR VPWR tag_array.tag0\[0\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_176_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13584_ clknet_leaf_61_clk _02213_ VGND VGND VPWR VPWR data_array.data0\[9\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_10796_ net3215 net1044 net505 VGND VGND VPWR VPWR _02541_ sky130_fd_sc_hd__mux2_1
XFILLER_13_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_171_3648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12535_ clknet_leaf_140_clk _01229_ VGND VGND VPWR VPWR tag_array.tag1\[11\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_129_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_916 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12466_ clknet_leaf_45_clk _01160_ VGND VGND VPWR VPWR data_array.data1\[9\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_132_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14205_ clknet_leaf_2_clk _02834_ VGND VGND VPWR VPWR data_array.data0\[2\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
X_11417_ clknet_leaf_270_clk _00227_ VGND VGND VPWR VPWR data_array.data0\[0\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_12397_ clknet_leaf_63_clk _01091_ VGND VGND VPWR VPWR data_array.data0\[14\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_153_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14136_ clknet_leaf_56_clk _02765_ VGND VGND VPWR VPWR data_array.data0\[1\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
X_11348_ net900 net4023 net798 VGND VGND VPWR VPWR _03091_ sky130_fd_sc_hd__mux2_1
X_14067_ clknet_leaf_44_clk _02696_ VGND VGND VPWR VPWR data_array.data1\[6\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
X_11279_ net914 net3455 net680 VGND VGND VPWR VPWR _03022_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13018_ clknet_leaf_89_clk _01712_ VGND VGND VPWR VPWR data_array.data0\[3\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_33_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05840_ net851 data_array.rdata0\[3\] net1148 VGND VGND VPWR VPWR _03354_ sky130_fd_sc_hd__o21a_1
XFILLER_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05771_ _03286_ _03287_ _03238_ _03269_ VGND VGND VPWR VPWR _03288_ sky130_fd_sc_hd__a211o_1
XFILLER_63_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07510_ data_array.data1\[0\]\[6\] net1329 net1235 data_array.data1\[3\]\[6\] _04744_
+ VGND VGND VPWR VPWR _04745_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_18_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08490_ net1718 net629 VGND VGND VPWR VPWR _00292_ sky130_fd_sc_hd__nand2b_1
XFILLER_23_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07441_ data_array.data1\[13\]\[0\] net1556 net1460 data_array.data1\[14\]\[0\] VGND
+ VGND VPWR VPWR _04682_ sky130_fd_sc_hd__a22o_1
X_07372_ net1193 _04613_ _04617_ net1619 VGND VGND VPWR VPWR _04620_ sky130_fd_sc_hd__a22o_1
XFILLER_128_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09111_ net1099 net4024 net568 VGND VGND VPWR VPWR _00865_ sky130_fd_sc_hd__mux2_1
X_06323_ tag_array.tag0\[13\]\[12\] net1597 net1501 tag_array.tag0\[14\]\[12\] VGND
+ VGND VPWR VPWR _03666_ sky130_fd_sc_hd__a22o_1
XFILLER_31_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09042_ net2020 net856 net421 VGND VGND VPWR VPWR _00797_ sky130_fd_sc_hd__mux2_1
XFILLER_108_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06254_ tag_array.tag0\[12\]\[6\] net1373 net1279 tag_array.tag0\[15\]\[6\] _03602_
+ VGND VGND VPWR VPWR _03603_ sky130_fd_sc_hd__a221o_1
XFILLER_159_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold400 data_array.data1\[0\]\[56\] VGND VGND VPWR VPWR net2051 sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 data_array.data1\[8\]\[41\] VGND VGND VPWR VPWR net2062 sky130_fd_sc_hd__dlygate4sd3_1
X_06185_ net1221 _03535_ _03539_ net1172 VGND VGND VPWR VPWR _03541_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_92_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold422 data_array.data1\[8\]\[61\] VGND VGND VPWR VPWR net2073 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold433 tag_array.tag0\[13\]\[21\] VGND VGND VPWR VPWR net2084 sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 data_array.data1\[1\]\[38\] VGND VGND VPWR VPWR net2095 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold455 tag_array.tag0\[10\]\[12\] VGND VGND VPWR VPWR net2106 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold466 data_array.data1\[1\]\[12\] VGND VGND VPWR VPWR net2117 sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 data_array.data0\[1\]\[34\] VGND VGND VPWR VPWR net2128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold488 data_array.data1\[4\]\[60\] VGND VGND VPWR VPWR net2139 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout902 _05524_ VGND VGND VPWR VPWR net902 sky130_fd_sc_hd__clkbuf_2
X_09944_ net1052 net3946 net376 VGND VGND VPWR VPWR _01693_ sky130_fd_sc_hd__mux2_1
XFILLER_131_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold499 data_array.data0\[8\]\[17\] VGND VGND VPWR VPWR net2150 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout913 _05518_ VGND VGND VPWR VPWR net913 sky130_fd_sc_hd__buf_1
Xfanout924 _05512_ VGND VGND VPWR VPWR net924 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_70_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout935 _05508_ VGND VGND VPWR VPWR net935 sky130_fd_sc_hd__buf_1
XFILLER_48_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout946 net947 VGND VGND VPWR VPWR net946 sky130_fd_sc_hd__clkbuf_2
XFILLER_38_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout957 net959 VGND VGND VPWR VPWR net957 sky130_fd_sc_hd__clkbuf_2
X_09875_ net970 net3035 net378 VGND VGND VPWR VPWR _01625_ sky130_fd_sc_hd__mux2_1
XFILLER_131_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout968 _05490_ VGND VGND VPWR VPWR net968 sky130_fd_sc_hd__clkbuf_2
Xhold1100 data_array.data0\[2\]\[38\] VGND VGND VPWR VPWR net2751 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout979 _05486_ VGND VGND VPWR VPWR net979 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1111 tag_array.tag0\[12\]\[8\] VGND VGND VPWR VPWR net2762 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1122 data_array.data1\[13\]\[4\] VGND VGND VPWR VPWR net2773 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_86_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08826_ net1950 net940 net448 VGND VGND VPWR VPWR _00584_ sky130_fd_sc_hd__mux2_1
Xhold1133 data_array.data1\[14\]\[14\] VGND VGND VPWR VPWR net2784 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_161_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1144 data_array.data0\[9\]\[12\] VGND VGND VPWR VPWR net2795 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1155 tag_array.tag0\[3\]\[6\] VGND VGND VPWR VPWR net2806 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1166 data_array.data1\[14\]\[49\] VGND VGND VPWR VPWR net2817 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1177 tag_array.tag1\[1\]\[24\] VGND VGND VPWR VPWR net2828 sky130_fd_sc_hd__dlygate4sd3_1
X_08757_ net695 net3142 net458 VGND VGND VPWR VPWR _00516_ sky130_fd_sc_hd__mux2_1
Xhold1188 data_array.data1\[2\]\[25\] VGND VGND VPWR VPWR net2839 sky130_fd_sc_hd__dlygate4sd3_1
X_05969_ data_array.rdata0\[46\] net846 net1143 VGND VGND VPWR VPWR _03440_ sky130_fd_sc_hd__o21a_1
Xhold1199 data_array.data0\[12\]\[47\] VGND VGND VPWR VPWR net2850 sky130_fd_sc_hd__dlygate4sd3_1
X_07708_ data_array.data1\[4\]\[24\] net1387 net1293 data_array.data1\[7\]\[24\] _04924_
+ VGND VGND VPWR VPWR _04925_ sky130_fd_sc_hd__a221o_1
X_08688_ net1824 net772 net487 VGND VGND VPWR VPWR _00447_ sky130_fd_sc_hd__mux2_1
XFILLER_54_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07639_ data_array.data1\[9\]\[18\] net1536 net1440 data_array.data1\[10\]\[18\]
+ VGND VGND VPWR VPWR _04862_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_105_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_170 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10650_ net2247 net862 net475 VGND VGND VPWR VPWR _02395_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_153_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1013 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09309_ net743 net2796 net546 VGND VGND VPWR VPWR _01063_ sky130_fd_sc_hd__mux2_1
X_10581_ net883 net4334 net454 VGND VGND VPWR VPWR _02326_ sky130_fd_sc_hd__mux2_1
X_12320_ clknet_leaf_252_clk _00022_ VGND VGND VPWR VPWR data_array.rdata0\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_182_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12251_ clknet_leaf_137_clk _01009_ VGND VGND VPWR VPWR tag_array.tag1\[14\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_181_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11202_ net966 net3925 net656 VGND VGND VPWR VPWR _02945_ sky130_fd_sc_hd__mux2_1
XFILLER_163_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12182_ clknet_leaf_169_clk _00990_ VGND VGND VPWR VPWR tag_array.tag0\[14\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_123_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11133_ net985 net2502 net548 VGND VGND VPWR VPWR _02876_ sky130_fd_sc_hd__mux2_1
XFILLER_122_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11064_ net1857 net1007 net331 VGND VGND VPWR VPWR _02807_ sky130_fd_sc_hd__mux2_1
XFILLER_49_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10015_ net1024 net3491 net555 VGND VGND VPWR VPWR _01764_ sky130_fd_sc_hd__mux2_1
XFILLER_48_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2390 data_array.data1\[11\]\[61\] VGND VGND VPWR VPWR net4041 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_92_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_125_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11966_ clknet_leaf_127_clk _00774_ VGND VGND VPWR VPWR data_array.data0\[4\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
X_13705_ clknet_leaf_267_clk _02334_ VGND VGND VPWR VPWR data_array.data1\[1\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_10917_ net1074 net3333 net532 VGND VGND VPWR VPWR _02662_ sky130_fd_sc_hd__mux2_1
X_11897_ clknet_leaf_243_clk _00705_ VGND VGND VPWR VPWR data_array.data0\[5\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_44_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13636_ clknet_leaf_206_clk _02265_ VGND VGND VPWR VPWR data_array.data0\[9\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
X_10848_ net1094 net3185 net520 VGND VGND VPWR VPWR _02593_ sky130_fd_sc_hd__mux2_1
XFILLER_158_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13567_ clknet_leaf_28_clk _02196_ VGND VGND VPWR VPWR tag_array.dirty1\[7\] sky130_fd_sc_hd__dfxtp_1
X_10779_ net858 net2536 net493 VGND VGND VPWR VPWR _02524_ sky130_fd_sc_hd__mux2_1
XFILLER_173_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Left_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12518_ clknet_leaf_95_clk _01212_ VGND VGND VPWR VPWR tag_array.tag1\[11\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_13498_ clknet_leaf_31_clk _02127_ VGND VGND VPWR VPWR tag_array.dirty1\[12\] sky130_fd_sc_hd__dfxtp_1
X_12449_ clknet_leaf_265_clk _01143_ VGND VGND VPWR VPWR data_array.data1\[9\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_154_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14119_ clknet_leaf_37_clk _02748_ VGND VGND VPWR VPWR data_array.data0\[1\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_07990_ _05180_ _05181_ VGND VGND VPWR VPWR _00107_ sky130_fd_sc_hd__or2_1
X_06941_ data_array.data0\[1\]\[18\] net1536 net1440 data_array.data0\[2\]\[18\] VGND
+ VGND VPWR VPWR _04228_ sky130_fd_sc_hd__a22o_1
XFILLER_119_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09660_ net749 net3164 net612 VGND VGND VPWR VPWR _01412_ sky130_fd_sc_hd__mux2_1
XFILLER_28_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06872_ data_array.data0\[0\]\[12\] net1386 net1292 data_array.data0\[3\]\[12\] _04164_
+ VGND VGND VPWR VPWR _04165_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_2_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08611_ net778 net4056 net517 VGND VGND VPWR VPWR _00370_ sky130_fd_sc_hd__mux2_1
XFILLER_95_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05823_ _03280_ _03282_ _03301_ _03312_ VGND VGND VPWR VPWR _03340_ sky130_fd_sc_hd__or4_1
X_09591_ net987 net3968 net398 VGND VGND VPWR VPWR _01343_ sky130_fd_sc_hd__mux2_1
X_08542_ net786 net4439 net580 VGND VGND VPWR VPWR _00310_ sky130_fd_sc_hd__mux2_1
X_05754_ net8 fsm.tag_out1\[9\] VGND VGND VPWR VPWR _03271_ sky130_fd_sc_hd__and2b_1
XFILLER_36_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_1043 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08473_ net1625 net1275 net814 net1701 VGND VGND VPWR VPWR _00287_ sky130_fd_sc_hd__a31o_1
X_05685_ _03198_ _03199_ _03200_ _03201_ VGND VGND VPWR VPWR _03202_ sky130_fd_sc_hd__or4_1
XFILLER_51_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07424_ data_array.data0\[12\]\[62\] net1412 net1318 data_array.data0\[15\]\[62\]
+ _04666_ VGND VGND VPWR VPWR _04667_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_46_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07355_ data_array.data0\[5\]\[56\] net1531 net1435 data_array.data0\[6\]\[56\] VGND
+ VGND VPWR VPWR _04604_ sky130_fd_sc_hd__a22o_1
XFILLER_137_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06306_ net1183 _03645_ _03649_ net1231 VGND VGND VPWR VPWR _03651_ sky130_fd_sc_hd__a22o_1
XFILLER_108_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07286_ _04540_ _04541_ VGND VGND VPWR VPWR _00043_ sky130_fd_sc_hd__or2_1
XFILLER_163_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09025_ net1893 net927 net418 VGND VGND VPWR VPWR _00780_ sky130_fd_sc_hd__mux2_1
XFILLER_108_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06237_ tag_array.tag0\[1\]\[4\] net1561 net1465 tag_array.tag0\[2\]\[4\] VGND VGND
+ VPWR VPWR _03588_ sky130_fd_sc_hd__a22o_1
XFILLER_152_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold230 data_array.data0\[0\]\[46\] VGND VGND VPWR VPWR net1881 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06168_ tag_array.valid0\[12\] net1408 net1314 tag_array.valid0\[15\] _03524_ VGND
+ VGND VPWR VPWR _03525_ sky130_fd_sc_hd__a221o_1
Xhold241 tag_array.tag1\[4\]\[21\] VGND VGND VPWR VPWR net1892 sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 data_array.data1\[1\]\[4\] VGND VGND VPWR VPWR net1903 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold263 data_array.data1\[2\]\[30\] VGND VGND VPWR VPWR net1914 sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 data_array.data0\[0\]\[8\] VGND VGND VPWR VPWR net1925 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold285 data_array.data1\[4\]\[0\] VGND VGND VPWR VPWR net1936 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_160_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold296 data_array.data1\[2\]\[39\] VGND VGND VPWR VPWR net1947 sky130_fd_sc_hd__dlygate4sd3_1
X_06099_ data_array.rdata0\[14\] net1140 net1114 data_array.rdata1\[14\] VGND VGND
+ VPWR VPWR net268 sky130_fd_sc_hd__a22o_1
XFILLER_172_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout710 net711 VGND VGND VPWR VPWR net710 sky130_fd_sc_hd__clkbuf_2
Xfanout721 _05401_ VGND VGND VPWR VPWR net721 sky130_fd_sc_hd__clkbuf_2
XFILLER_49_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout732 _05395_ VGND VGND VPWR VPWR net732 sky130_fd_sc_hd__clkbuf_2
X_09927_ net698 net2124 net603 VGND VGND VPWR VPWR _01677_ sky130_fd_sc_hd__mux2_1
Xfanout743 _05389_ VGND VGND VPWR VPWR net743 sky130_fd_sc_hd__buf_1
Xfanout754 net755 VGND VGND VPWR VPWR net754 sky130_fd_sc_hd__clkbuf_2
Xfanout765 _05379_ VGND VGND VPWR VPWR net765 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_146_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout776 _05373_ VGND VGND VPWR VPWR net776 sky130_fd_sc_hd__clkbuf_2
XFILLER_74_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09858_ net1037 net3659 net379 VGND VGND VPWR VPWR _01608_ sky130_fd_sc_hd__mux2_1
Xfanout787 net788 VGND VGND VPWR VPWR net787 sky130_fd_sc_hd__buf_1
XFILLER_105_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout798 net799 VGND VGND VPWR VPWR net798 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_107_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08809_ net2049 net1009 net442 VGND VGND VPWR VPWR _00567_ sky130_fd_sc_hd__mux2_1
X_09789_ net1053 net4032 net390 VGND VGND VPWR VPWR _01540_ sky130_fd_sc_hd__mux2_1
XFILLER_22_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11820_ clknet_leaf_8_clk _00628_ VGND VGND VPWR VPWR data_array.data0\[7\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_11751_ clknet_leaf_249_clk _00559_ VGND VGND VPWR VPWR data_array.data0\[8\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_80_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_80_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_81_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10702_ net2350 net908 net480 VGND VGND VPWR VPWR _02447_ sky130_fd_sc_hd__mux2_1
XFILLER_14_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14470_ clknet_leaf_215_clk _03093_ VGND VGND VPWR VPWR data_array.data1\[7\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_120_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11682_ clknet_leaf_128_clk _00490_ VGND VGND VPWR VPWR tag_array.tag1\[1\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_41_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13421_ clknet_leaf_259_clk _02051_ VGND VGND VPWR VPWR data_array.data1\[8\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
X_10633_ net1956 net930 net467 VGND VGND VPWR VPWR _02378_ sky130_fd_sc_hd__mux2_1
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13352_ clknet_leaf_206_clk _01982_ VGND VGND VPWR VPWR data_array.data0\[10\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
X_10564_ net950 net4331 net463 VGND VGND VPWR VPWR _02309_ sky130_fd_sc_hd__mux2_1
XFILLER_128_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12303_ clknet_leaf_105_clk _01061_ VGND VGND VPWR VPWR tag_array.tag1\[12\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_20_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13283_ clknet_leaf_9_clk _01913_ VGND VGND VPWR VPWR data_array.data0\[11\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
X_10495_ net965 net3432 net350 VGND VGND VPWR VPWR _02240_ sky130_fd_sc_hd__mux2_1
X_12234_ clknet_leaf_147_clk _00163_ VGND VGND VPWR VPWR fsm.tag_out1\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_122_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12165_ clknet_leaf_182_clk _00973_ VGND VGND VPWR VPWR tag_array.tag0\[13\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_166_3547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11116_ net1054 net2866 net548 VGND VGND VPWR VPWR _02859_ sky130_fd_sc_hd__mux2_1
X_12096_ clknet_leaf_84_clk _00904_ VGND VGND VPWR VPWR data_array.data1\[14\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_49_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_183_3872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_890 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_3883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_127_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11047_ net1791 net1072 net333 VGND VGND VPWR VPWR _02790_ sky130_fd_sc_hd__mux2_1
XFILLER_37_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput9 cpu_addr[17] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_4
XFILLER_49_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12998_ clknet_leaf_225_clk _01692_ VGND VGND VPWR VPWR data_array.data0\[3\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_45_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11949_ clknet_leaf_176_clk _00757_ VGND VGND VPWR VPWR data_array.data0\[4\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_71_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_71_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_44_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13619_ clknet_leaf_84_clk _02248_ VGND VGND VPWR VPWR data_array.data0\[9\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07140_ data_array.data0\[0\]\[36\] net1413 net1319 data_array.data0\[3\]\[36\] _04408_
+ VGND VGND VPWR VPWR _04409_ sky130_fd_sc_hd__a221o_1
XFILLER_125_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_735 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07071_ data_array.data0\[13\]\[30\] net1581 net1485 data_array.data0\[14\]\[30\]
+ VGND VGND VPWR VPWR _04346_ sky130_fd_sc_hd__a22o_1
X_06022_ net158 net1153 _03474_ _03475_ VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__a22o_1
Xoutput302 net302 VGND VGND VPWR VPWR mem_wdata[45] sky130_fd_sc_hd__buf_2
Xoutput313 net313 VGND VGND VPWR VPWR mem_wdata[55] sky130_fd_sc_hd__buf_2
Xoutput324 net324 VGND VGND VPWR VPWR mem_wdata[7] sky130_fd_sc_hd__buf_2
XFILLER_154_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07973_ data_array.data1\[13\]\[48\] net1590 net1494 data_array.data1\[14\]\[48\]
+ VGND VGND VPWR VPWR _05166_ sky130_fd_sc_hd__a22o_1
X_09712_ net738 net3548 net610 VGND VGND VPWR VPWR _01464_ sky130_fd_sc_hd__mux2_1
X_06924_ data_array.data0\[13\]\[17\] net1528 net1432 data_array.data0\[14\]\[17\]
+ VGND VGND VPWR VPWR _04212_ sky130_fd_sc_hd__a22o_1
XFILLER_110_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09643_ net716 net3720 net616 VGND VGND VPWR VPWR _01395_ sky130_fd_sc_hd__mux2_1
X_06855_ net1635 _04143_ _04147_ net1209 VGND VGND VPWR VPWR _04150_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_48_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05806_ net24 fsm.tag_out0\[23\] VGND VGND VPWR VPWR _03323_ sky130_fd_sc_hd__and2b_1
X_09574_ net1052 net4446 net398 VGND VGND VPWR VPWR _01326_ sky130_fd_sc_hd__mux2_1
X_06786_ data_array.data0\[12\]\[4\] net1391 net1297 data_array.data0\[15\]\[4\] _04086_
+ VGND VGND VPWR VPWR _04087_ sky130_fd_sc_hd__a221o_1
XFILLER_70_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08525_ _03509_ _03519_ net821 VGND VGND VPWR VPWR _05588_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_65_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05737_ _03143_ fsm.tag_out1\[20\] _03247_ _03248_ _03253_ VGND VGND VPWR VPWR _03254_
+ sky130_fd_sc_hd__a2111o_1
XFILLER_36_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_62_clk clknet_5_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_62_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_168_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08456_ net1992 net868 net693 VGND VGND VPWR VPWR _00281_ sky130_fd_sc_hd__mux2_1
XFILLER_24_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_05668_ net10 fsm.tag_out0\[11\] VGND VGND VPWR VPWR _03185_ sky130_fd_sc_hd__and2b_1
XFILLER_51_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07407_ _04650_ _04651_ VGND VGND VPWR VPWR _00056_ sky130_fd_sc_hd__or2_1
XFILLER_51_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08387_ net2742 net962 net688 VGND VGND VPWR VPWR _00258_ sky130_fd_sc_hd__mux2_1
XFILLER_183_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_871 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07338_ data_array.data0\[4\]\[54\] net1356 net1262 data_array.data0\[7\]\[54\] _04588_
+ VGND VGND VPWR VPWR _04589_ sky130_fd_sc_hd__a221o_1
XFILLER_136_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07269_ data_array.data0\[13\]\[48\] net1581 net1485 data_array.data0\[14\]\[48\]
+ VGND VGND VPWR VPWR _04526_ sky130_fd_sc_hd__a22o_1
X_09008_ net2256 net992 net422 VGND VGND VPWR VPWR _00763_ sky130_fd_sc_hd__mux2_1
XFILLER_3_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10280_ net2158 net1041 net634 VGND VGND VPWR VPWR _02027_ sky130_fd_sc_hd__mux2_1
XFILLER_117_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_148_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1505 net1507 VGND VGND VPWR VPWR net1505 sky130_fd_sc_hd__clkbuf_4
Xfanout1516 net1517 VGND VGND VPWR VPWR net1516 sky130_fd_sc_hd__buf_2
Xfanout1527 net1529 VGND VGND VPWR VPWR net1527 sky130_fd_sc_hd__clkbuf_4
Xfanout1538 net1539 VGND VGND VPWR VPWR net1538 sky130_fd_sc_hd__clkbuf_4
Xfanout540 _05597_ VGND VGND VPWR VPWR net540 sky130_fd_sc_hd__buf_4
XFILLER_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout551 net552 VGND VGND VPWR VPWR net551 sky130_fd_sc_hd__buf_4
XFILLER_116_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1549 net1554 VGND VGND VPWR VPWR net1549 sky130_fd_sc_hd__buf_2
Xfanout562 net563 VGND VGND VPWR VPWR net562 sky130_fd_sc_hd__buf_4
X_13970_ clknet_leaf_116_clk _02599_ VGND VGND VPWR VPWR data_array.data1\[5\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout573 net575 VGND VGND VPWR VPWR net573 sky130_fd_sc_hd__clkbuf_8
XFILLER_120_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout584 _05591_ VGND VGND VPWR VPWR net584 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_161_3455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout595 net598 VGND VGND VPWR VPWR net595 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_161_3466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12921_ clknet_leaf_262_clk _01615_ VGND VGND VPWR VPWR data_array.data0\[13\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ clknet_leaf_128_clk _01546_ VGND VGND VPWR VPWR data_array.data0\[12\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_55_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11803_ clknet_leaf_210_clk _00611_ VGND VGND VPWR VPWR data_array.data0\[7\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_73_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12783_ clknet_leaf_233_clk _01477_ VGND VGND VPWR VPWR tag_array.tag1\[10\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_53_clk clknet_5_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_53_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_42_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11734_ clknet_leaf_227_clk _00542_ VGND VGND VPWR VPWR data_array.data0\[8\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14453_ clknet_leaf_217_clk _03076_ VGND VGND VPWR VPWR data_array.data1\[7\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
X_11665_ clknet_leaf_195_clk _00473_ VGND VGND VPWR VPWR tag_array.tag1\[1\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_175_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_6_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_6_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_30_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10616_ net2625 net997 net467 VGND VGND VPWR VPWR _02361_ sky130_fd_sc_hd__mux2_1
XFILLER_128_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13404_ clknet_leaf_88_clk _02034_ VGND VGND VPWR VPWR data_array.data1\[8\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14384_ clknet_leaf_6_clk _03007_ VGND VGND VPWR VPWR data_array.data1\[10\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
X_11596_ clknet_leaf_166_clk _00404_ VGND VGND VPWR VPWR tag_array.tag1\[4\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13335_ clknet_leaf_84_clk _01965_ VGND VGND VPWR VPWR data_array.data0\[10\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10547_ net1016 net2362 net457 VGND VGND VPWR VPWR _02292_ sky130_fd_sc_hd__mux2_1
XFILLER_41_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13266_ clknet_leaf_235_clk _01896_ VGND VGND VPWR VPWR data_array.data0\[11\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_94_Left_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10478_ net1032 net4568 net349 VGND VGND VPWR VPWR _02223_ sky130_fd_sc_hd__mux2_1
XFILLER_136_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12217_ clknet_leaf_184_clk _00147_ VGND VGND VPWR VPWR fsm.tag_out0\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_124_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13197_ clknet_leaf_11_clk _00091_ VGND VGND VPWR VPWR data_array.rdata1\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_68_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12148_ clknet_leaf_144_clk _00956_ VGND VGND VPWR VPWR tag_array.tag0\[13\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_155_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12079_ clknet_leaf_263_clk _00887_ VGND VGND VPWR VPWR data_array.data1\[14\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_139_Right_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06640_ tag_array.tag1\[1\]\[16\] net1609 net1513 tag_array.tag1\[2\]\[16\] VGND
+ VGND VPWR VPWR _03954_ sky130_fd_sc_hd__a22o_1
XFILLER_37_479 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06571_ _03890_ _03891_ VGND VGND VPWR VPWR _00180_ sky130_fd_sc_hd__or2_1
XFILLER_75_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_44_clk clknet_5_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_44_clk sky130_fd_sc_hd__clkbuf_8
X_08310_ net102 net37 net1641 VGND VGND VPWR VPWR _05443_ sky130_fd_sc_hd__mux2_1
XFILLER_75_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09290_ net718 net2637 net559 VGND VGND VPWR VPWR _01044_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08241_ net730 net4156 net803 VGND VGND VPWR VPWR _00211_ sky130_fd_sc_hd__mux2_1
XANTENNA_14 _03132_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_25 _05399_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_36 net390 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_47 net659 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_58 net1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08172_ lru_array.lru_mem\[8\] net1373 net1279 lru_array.lru_mem\[11\] _05346_ VGND
+ VGND VPWR VPWR _05347_ sky130_fd_sc_hd__a221o_1
XFILLER_119_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_69 _00022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07123_ data_array.data0\[12\]\[35\] net1346 net1252 data_array.data0\[15\]\[35\]
+ _04392_ VGND VGND VPWR VPWR _04393_ sky130_fd_sc_hd__a221o_1
XFILLER_118_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07054_ net1169 _04325_ _04329_ net1217 VGND VGND VPWR VPWR _04331_ sky130_fd_sc_hd__a22o_1
X_06005_ data_array.rdata0\[58\] net849 net1144 VGND VGND VPWR VPWR _03464_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_58_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput165 net165 VGND VGND VPWR VPWR cpu_rdata[0] sky130_fd_sc_hd__buf_2
XFILLER_0_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput176 net176 VGND VGND VPWR VPWR cpu_rdata[1] sky130_fd_sc_hd__buf_4
XFILLER_114_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput187 net187 VGND VGND VPWR VPWR cpu_rdata[2] sky130_fd_sc_hd__clkbuf_4
Xhold2901 data_array.data1\[15\]\[35\] VGND VGND VPWR VPWR net4552 sky130_fd_sc_hd__dlygate4sd3_1
Xoutput198 net198 VGND VGND VPWR VPWR cpu_rdata[3] sky130_fd_sc_hd__buf_6
Xhold2912 tag_array.tag0\[10\]\[19\] VGND VGND VPWR VPWR net4563 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_141_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2923 data_array.data0\[9\]\[63\] VGND VGND VPWR VPWR net4574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2934 tag_array.tag1\[10\]\[3\] VGND VGND VPWR VPWR net4585 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2945 data_array.data1\[10\]\[29\] VGND VGND VPWR VPWR net4596 sky130_fd_sc_hd__dlygate4sd3_1
X_07956_ net1165 _05145_ _05149_ net1213 VGND VGND VPWR VPWR _05151_ sky130_fd_sc_hd__a22o_1
Xhold2956 data_array.data0\[5\]\[54\] VGND VGND VPWR VPWR net4607 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2967 data_array.data0\[14\]\[45\] VGND VGND VPWR VPWR net4618 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_101_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06907_ data_array.data0\[12\]\[15\] net1390 net1296 data_array.data0\[15\]\[15\]
+ _04196_ VGND VGND VPWR VPWR _04197_ sky130_fd_sc_hd__a221o_1
XFILLER_46_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_733 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07887_ data_array.data1\[1\]\[40\] net1606 net1510 data_array.data1\[2\]\[40\] VGND
+ VGND VPWR VPWR _05088_ sky130_fd_sc_hd__a22o_1
XFILLER_28_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_106_Right_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06838_ data_array.data0\[5\]\[9\] net1580 net1484 data_array.data0\[6\]\[9\] VGND
+ VGND VPWR VPWR _04134_ sky130_fd_sc_hd__a22o_1
X_09626_ net784 net3374 net615 VGND VGND VPWR VPWR _01378_ sky130_fd_sc_hd__mux2_1
XFILLER_44_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09557_ net699 net4327 net619 VGND VGND VPWR VPWR _01310_ sky130_fd_sc_hd__mux2_1
X_06769_ _04070_ _04071_ VGND VGND VPWR VPWR _00022_ sky130_fd_sc_hd__or2_1
XFILLER_71_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_35_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_8
X_08508_ net821 net811 net854 _05574_ VGND VGND VPWR VPWR _05576_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_80_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09488_ net776 net2814 net624 VGND VGND VPWR VPWR _01241_ sky130_fd_sc_hd__mux2_1
XFILLER_12_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08439_ net149 net84 net1639 VGND VGND VPWR VPWR _05529_ sky130_fd_sc_hd__mux2_1
XFILLER_156_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11450_ clknet_leaf_236_clk _00260_ VGND VGND VPWR VPWR data_array.data0\[0\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10401_ net1735 net1050 net668 VGND VGND VPWR VPWR _02147_ sky130_fd_sc_hd__mux2_1
X_11381_ net164 VGND VGND VPWR VPWR _00191_ sky130_fd_sc_hd__inv_2
XFILLER_180_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13120_ clknet_leaf_142_clk _01814_ VGND VGND VPWR VPWR tag_array.tag0\[3\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_10332_ net770 net4181 net592 VGND VGND VPWR VPWR _02079_ sky130_fd_sc_hd__mux2_1
XFILLER_180_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13051_ clknet_leaf_251_clk _01745_ VGND VGND VPWR VPWR data_array.data1\[13\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_10263_ net3598 net1111 net638 VGND VGND VPWR VPWR _02010_ sky130_fd_sc_hd__mux2_1
XFILLER_152_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12002_ clknet_leaf_95_clk _00810_ VGND VGND VPWR VPWR data_array.data0\[6\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_127_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1302 net1305 VGND VGND VPWR VPWR net1302 sky130_fd_sc_hd__clkbuf_4
X_10194_ net1029 net2934 net360 VGND VGND VPWR VPWR _01941_ sky130_fd_sc_hd__mux2_1
XFILLER_78_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1313 net1314 VGND VGND VPWR VPWR net1313 sky130_fd_sc_hd__clkbuf_4
Xfanout1324 net1327 VGND VGND VPWR VPWR net1324 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_180_3820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1335 net1336 VGND VGND VPWR VPWR net1335 sky130_fd_sc_hd__clkbuf_4
Xfanout1346 net1348 VGND VGND VPWR VPWR net1346 sky130_fd_sc_hd__clkbuf_4
Xfanout1357 net1358 VGND VGND VPWR VPWR net1357 sky130_fd_sc_hd__clkbuf_4
Xfanout370 net374 VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__buf_4
XFILLER_47_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1368 net1370 VGND VGND VPWR VPWR net1368 sky130_fd_sc_hd__clkbuf_4
XFILLER_87_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout381 net385 VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__buf_4
Xfanout1379 net1382 VGND VGND VPWR VPWR net1379 sky130_fd_sc_hd__clkbuf_4
XFILLER_143_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout392 net393 VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__clkbuf_8
X_13953_ clknet_leaf_249_clk _02582_ VGND VGND VPWR VPWR data_array.data1\[4\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_93_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12904_ clknet_leaf_18_clk _01598_ VGND VGND VPWR VPWR data_array.data0\[13\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_13884_ clknet_leaf_212_clk _02513_ VGND VGND VPWR VPWR data_array.data1\[3\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12835_ clknet_leaf_46_clk _01529_ VGND VGND VPWR VPWR data_array.data0\[12\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_26_clk clknet_5_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_178_3771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_3782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ clknet_leaf_160_clk _01460_ VGND VGND VPWR VPWR tag_array.tag0\[6\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11717_ clknet_leaf_137_clk _00525_ VGND VGND VPWR VPWR tag_array.tag0\[9\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_12697_ clknet_leaf_162_clk _01391_ VGND VGND VPWR VPWR tag_array.tag0\[8\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_147_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14436_ clknet_leaf_130_clk _03059_ VGND VGND VPWR VPWR data_array.data1\[7\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_11648_ clknet_leaf_168_clk _00456_ VGND VGND VPWR VPWR tag_array.tag1\[2\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput12 cpu_addr[1] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
Xinput23 cpu_addr[2] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_1
Xinput34 cpu_wdata[0] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_1
Xinput45 cpu_wdata[1] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_1
X_14367_ clknet_leaf_254_clk _02990_ VGND VGND VPWR VPWR data_array.data1\[10\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_11579_ clknet_leaf_234_clk _00387_ VGND VGND VPWR VPWR tag_array.tag1\[5\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_155_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput56 cpu_wdata[2] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_1
XFILLER_155_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold807 data_array.data1\[15\]\[54\] VGND VGND VPWR VPWR net2458 sky130_fd_sc_hd__dlygate4sd3_1
Xinput67 cpu_wdata[3] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_1
Xinput78 cpu_wdata[4] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_1
Xinput89 cpu_wdata[5] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__clkbuf_1
X_13318_ clknet_leaf_229_clk _01948_ VGND VGND VPWR VPWR data_array.data0\[10\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold818 data_array.data0\[12\]\[12\] VGND VGND VPWR VPWR net2469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold829 data_array.data0\[6\]\[28\] VGND VGND VPWR VPWR net2480 sky130_fd_sc_hd__dlygate4sd3_1
X_14298_ clknet_leaf_19_clk _02927_ VGND VGND VPWR VPWR data_array.data1\[11\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_182_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13249_ clknet_leaf_22_clk _01879_ VGND VGND VPWR VPWR data_array.data0\[11\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_69_302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2208 data_array.data1\[3\]\[61\] VGND VGND VPWR VPWR net3859 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2219 data_array.data1\[8\]\[57\] VGND VGND VPWR VPWR net3870 sky130_fd_sc_hd__dlygate4sd3_1
X_07810_ data_array.data1\[5\]\[33\] net1588 net1492 data_array.data1\[6\]\[33\] VGND
+ VGND VPWR VPWR _05018_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_36_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1507 data_array.data1\[9\]\[12\] VGND VGND VPWR VPWR net3158 sky130_fd_sc_hd__dlygate4sd3_1
X_08790_ net2268 net1087 net442 VGND VGND VPWR VPWR _00548_ sky130_fd_sc_hd__mux2_1
Xhold1518 tag_array.tag0\[5\]\[3\] VGND VGND VPWR VPWR net3169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1529 data_array.data0\[6\]\[63\] VGND VGND VPWR VPWR net3180 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_81_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07741_ data_array.data1\[0\]\[27\] net1356 net1262 data_array.data1\[3\]\[27\] _04954_
+ VGND VGND VPWR VPWR _04955_ sky130_fd_sc_hd__a221o_1
XFILLER_111_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07672_ data_array.data1\[9\]\[21\] net1547 net1451 data_array.data1\[10\]\[21\]
+ VGND VGND VPWR VPWR _04892_ sky130_fd_sc_hd__a22o_1
X_09411_ net1021 net3986 net580 VGND VGND VPWR VPWR _01164_ sky130_fd_sc_hd__mux2_1
XFILLER_16_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06623_ tag_array.tag1\[4\]\[14\] net1368 net1274 tag_array.tag1\[7\]\[14\] _03938_
+ VGND VGND VPWR VPWR _03939_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_17_clk clknet_5_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_8
X_09342_ net1033 net2462 net407 VGND VGND VPWR VPWR _01095_ sky130_fd_sc_hd__mux2_1
XFILLER_179_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06554_ tag_array.tag1\[13\]\[8\] net1608 net1512 tag_array.tag1\[14\]\[8\] VGND
+ VGND VPWR VPWR _03876_ sky130_fd_sc_hd__a22o_1
XFILLER_21_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09273_ net786 net3291 net556 VGND VGND VPWR VPWR _01027_ sky130_fd_sc_hd__mux2_1
X_06485_ tag_array.tag1\[8\]\[2\] net1388 net1294 tag_array.tag1\[11\]\[2\] _03812_
+ VGND VGND VPWR VPWR _03813_ sky130_fd_sc_hd__a221o_1
XFILLER_138_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08224_ net1650 net1161 net9 VGND VGND VPWR VPWR _05384_ sky130_fd_sc_hd__and3_1
XFILLER_178_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08155_ _05330_ _05331_ VGND VGND VPWR VPWR _00130_ sky130_fd_sc_hd__or2_1
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07106_ data_array.data0\[5\]\[33\] net1577 net1481 data_array.data0\[6\]\[33\] VGND
+ VGND VPWR VPWR _04378_ sky130_fd_sc_hd__a22o_1
X_08086_ data_array.data1\[0\]\[58\] net1359 net1265 data_array.data1\[3\]\[58\] _05268_
+ VGND VGND VPWR VPWR _05269_ sky130_fd_sc_hd__a221o_1
XFILLER_164_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07037_ data_array.data0\[0\]\[27\] net1347 net1253 data_array.data0\[3\]\[27\] _04314_
+ VGND VGND VPWR VPWR _04315_ sky130_fd_sc_hd__a221o_1
XFILLER_103_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2720 data_array.data0\[14\]\[35\] VGND VGND VPWR VPWR net4371 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_110_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2731 data_array.data1\[7\]\[51\] VGND VGND VPWR VPWR net4382 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2742 data_array.data1\[12\]\[29\] VGND VGND VPWR VPWR net4393 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_180_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08988_ net1809 net1072 net422 VGND VGND VPWR VPWR _00743_ sky130_fd_sc_hd__mux2_1
Xhold2753 data_array.data0\[10\]\[27\] VGND VGND VPWR VPWR net4404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2764 data_array.data1\[10\]\[34\] VGND VGND VPWR VPWR net4415 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2775 tag_array.tag0\[8\]\[7\] VGND VGND VPWR VPWR net4426 sky130_fd_sc_hd__dlygate4sd3_1
X_07939_ data_array.data1\[0\]\[45\] net1350 net1256 data_array.data1\[3\]\[45\] _05134_
+ VGND VGND VPWR VPWR _05135_ sky130_fd_sc_hd__a221o_1
Xhold2786 data_array.data0\[3\]\[55\] VGND VGND VPWR VPWR net4437 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2797 data_array.data1\[7\]\[3\] VGND VGND VPWR VPWR net4448 sky130_fd_sc_hd__dlygate4sd3_1
X_10950_ net942 net4291 net533 VGND VGND VPWR VPWR _02695_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_24 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09609_ net912 net4484 net399 VGND VGND VPWR VPWR _01361_ sky130_fd_sc_hd__mux2_1
X_10881_ net960 net3689 net516 VGND VGND VPWR VPWR _02626_ sky130_fd_sc_hd__mux2_1
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12620_ clknet_leaf_248_clk _01314_ VGND VGND VPWR VPWR data_array.data0\[15\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_43_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_159_Left_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_156_3354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12551_ clknet_leaf_147_clk _01245_ VGND VGND VPWR VPWR tag_array.tag0\[11\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_156_3365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11502_ clknet_leaf_233_clk _00310_ VGND VGND VPWR VPWR tag_array.tag1\[9\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_12482_ clknet_leaf_7_clk _01176_ VGND VGND VPWR VPWR data_array.data1\[9\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_117_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_997 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14221_ clknet_leaf_197_clk _02850_ VGND VGND VPWR VPWR data_array.data1\[12\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_11433_ clknet_leaf_8_clk _00243_ VGND VGND VPWR VPWR data_array.data0\[0\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14152_ clknet_leaf_230_clk _02781_ VGND VGND VPWR VPWR data_array.data0\[2\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_11364_ net1646 net4176 net600 VGND VGND VPWR VPWR _03107_ sky130_fd_sc_hd__mux2_1
XFILLER_125_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13103_ clknet_leaf_216_clk _01797_ VGND VGND VPWR VPWR data_array.data1\[13\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
X_10315_ net1831 net901 net637 VGND VGND VPWR VPWR _02062_ sky130_fd_sc_hd__mux2_1
X_14083_ clknet_leaf_54_clk _02712_ VGND VGND VPWR VPWR data_array.data1\[6\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
X_11295_ net820 net3102 _05553_ VGND VGND VPWR VPWR _03038_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_168_Left_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13034_ clknet_leaf_53_clk _01728_ VGND VGND VPWR VPWR data_array.data0\[3\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
X_10246_ net758 net3145 net597 VGND VGND VPWR VPWR _01993_ sky130_fd_sc_hd__mux2_1
XFILLER_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1110 _05420_ VGND VGND VPWR VPWR net1110 sky130_fd_sc_hd__clkbuf_2
XFILLER_78_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1121 net1122 VGND VGND VPWR VPWR net1121 sky130_fd_sc_hd__buf_2
Xfanout1132 net1133 VGND VGND VPWR VPWR net1132 sky130_fd_sc_hd__clkbuf_4
XFILLER_121_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10177_ net1096 net3218 net358 VGND VGND VPWR VPWR _01924_ sky130_fd_sc_hd__mux2_1
Xfanout1143 net1146 VGND VGND VPWR VPWR net1143 sky130_fd_sc_hd__buf_4
Xfanout1154 _03153_ VGND VGND VPWR VPWR net1154 sky130_fd_sc_hd__buf_8
XFILLER_120_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1165 net1167 VGND VGND VPWR VPWR net1165 sky130_fd_sc_hd__buf_4
Xfanout1176 net1177 VGND VGND VPWR VPWR net1176 sky130_fd_sc_hd__buf_4
Xfanout1187 _03526_ VGND VGND VPWR VPWR net1187 sky130_fd_sc_hd__buf_4
Xfanout1198 net1201 VGND VGND VPWR VPWR net1198 sky130_fd_sc_hd__buf_2
XFILLER_81_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13936_ clknet_leaf_123_clk _02565_ VGND VGND VPWR VPWR data_array.data1\[4\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_93_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13867_ clknet_leaf_256_clk _02496_ VGND VGND VPWR VPWR data_array.data1\[3\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_177_Left_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12818_ clknet_leaf_33_clk _01512_ VGND VGND VPWR VPWR tag_array.tag1\[0\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13798_ clknet_leaf_66_clk _02427_ VGND VGND VPWR VPWR data_array.data1\[2\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_12749_ clknet_leaf_109_clk _01443_ VGND VGND VPWR VPWR tag_array.tag0\[5\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_176_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06270_ tag_array.tag0\[5\]\[7\] net1607 net1511 tag_array.tag0\[6\]\[7\] VGND VGND
+ VPWR VPWR _03618_ sky130_fd_sc_hd__a22o_1
XFILLER_129_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14419_ clknet_leaf_28_clk _03042_ VGND VGND VPWR VPWR data_array.data1\[7\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold604 data_array.data0\[0\]\[56\] VGND VGND VPWR VPWR net2255 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold615 data_array.data0\[0\]\[3\] VGND VGND VPWR VPWR net2266 sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 data_array.data1\[1\]\[56\] VGND VGND VPWR VPWR net2277 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold637 data_array.data1\[8\]\[40\] VGND VGND VPWR VPWR net2288 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_94_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold648 data_array.data1\[4\]\[30\] VGND VGND VPWR VPWR net2299 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09960_ net988 net3223 net375 VGND VGND VPWR VPWR _01709_ sky130_fd_sc_hd__mux2_1
Xhold659 data_array.data0\[2\]\[3\] VGND VGND VPWR VPWR net2310 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_6_clk clknet_5_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_55_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08911_ net860 net3527 net441 VGND VGND VPWR VPWR _00668_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09891_ net905 net3856 net378 VGND VGND VPWR VPWR _01641_ sky130_fd_sc_hd__mux2_1
XFILLER_69_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_90_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2005 tag_array.tag0\[6\]\[19\] VGND VGND VPWR VPWR net3656 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2016 data_array.data0\[3\]\[17\] VGND VGND VPWR VPWR net3667 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2027 tag_array.tag0\[0\]\[12\] VGND VGND VPWR VPWR net3678 sky130_fd_sc_hd__dlygate4sd3_1
X_08842_ net3235 net876 net445 VGND VGND VPWR VPWR _00600_ sky130_fd_sc_hd__mux2_1
Xhold2038 data_array.data1\[5\]\[37\] VGND VGND VPWR VPWR net3689 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1304 data_array.data1\[7\]\[22\] VGND VGND VPWR VPWR net2955 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2049 tag_array.tag1\[5\]\[12\] VGND VGND VPWR VPWR net3700 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1315 data_array.data0\[5\]\[6\] VGND VGND VPWR VPWR net2966 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1326 data_array.data1\[13\]\[48\] VGND VGND VPWR VPWR net2977 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1337 data_array.data1\[9\]\[2\] VGND VGND VPWR VPWR net2988 sky130_fd_sc_hd__dlygate4sd3_1
X_08773_ net733 net3507 net451 VGND VGND VPWR VPWR _00532_ sky130_fd_sc_hd__mux2_1
Xhold1348 data_array.data0\[14\]\[60\] VGND VGND VPWR VPWR net2999 sky130_fd_sc_hd__dlygate4sd3_1
X_05985_ data_array.rdata1\[51\] net828 net837 VGND VGND VPWR VPWR _03451_ sky130_fd_sc_hd__a21o_1
Xhold1359 tag_array.tag0\[7\]\[9\] VGND VGND VPWR VPWR net3010 sky130_fd_sc_hd__dlygate4sd3_1
X_07724_ net1188 _04933_ _04937_ net1614 VGND VGND VPWR VPWR _04940_ sky130_fd_sc_hd__a22o_1
XFILLER_150_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07655_ data_array.data1\[8\]\[19\] net1394 net1300 data_array.data1\[11\]\[19\]
+ _04876_ VGND VGND VPWR VPWR _04877_ sky130_fd_sc_hd__a221o_1
XFILLER_25_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_864 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06606_ tag_array.tag1\[12\]\[13\] net1420 net1326 tag_array.tag1\[15\]\[13\] _03922_
+ VGND VGND VPWR VPWR _03923_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_0_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07586_ data_array.data1\[1\]\[13\] net1551 net1455 data_array.data1\[2\]\[13\] VGND
+ VGND VPWR VPWR _04814_ sky130_fd_sc_hd__a22o_1
XFILLER_80_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_16 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09325_ net1103 net3437 net404 VGND VGND VPWR VPWR _01078_ sky130_fd_sc_hd__mux2_1
X_06537_ net1219 _03855_ _03859_ net1172 VGND VGND VPWR VPWR _03861_ sky130_fd_sc_hd__a22o_1
XFILLER_167_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclone15 net851 VGND VGND VPWR VPWR net1666 sky130_fd_sc_hd__buf_6
XFILLER_167_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09256_ net756 net3811 net576 VGND VGND VPWR VPWR _01010_ sky130_fd_sc_hd__mux2_1
X_06468_ tag_array.tag1\[5\]\[0\] net1575 net1479 tag_array.tag1\[6\]\[0\] VGND VGND
+ VPWR VPWR _03798_ sky130_fd_sc_hd__a22o_1
X_08207_ fsm.tag_out1\[4\] net816 net808 fsm.tag_out0\[4\] _05372_ VGND VGND VPWR
+ VPWR _05373_ sky130_fd_sc_hd__a221o_2
XFILLER_182_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09187_ net732 net3186 net627 VGND VGND VPWR VPWR _00941_ sky130_fd_sc_hd__mux2_1
X_06399_ tag_array.tag0\[0\]\[19\] net1404 net1310 tag_array.tag0\[3\]\[19\] _03734_
+ VGND VGND VPWR VPWR _03735_ sky130_fd_sc_hd__a221o_1
XFILLER_175_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08138_ data_array.data1\[9\]\[63\] net1553 net1457 data_array.data1\[10\]\[63\]
+ VGND VGND VPWR VPWR _05316_ sky130_fd_sc_hd__a22o_1
XFILLER_175_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08069_ data_array.data1\[12\]\[57\] net1347 net1253 data_array.data1\[15\]\[57\]
+ _05252_ VGND VGND VPWR VPWR _05253_ sky130_fd_sc_hd__a221o_1
XFILLER_161_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10100_ net2214 net725 net642 VGND VGND VPWR VPWR _01849_ sky130_fd_sc_hd__mux2_1
XFILLER_134_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11080_ net1830 net940 net335 VGND VGND VPWR VPWR _02823_ sky130_fd_sc_hd__mux2_1
XFILLER_89_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10031_ net960 net3779 net554 VGND VGND VPWR VPWR _01780_ sky130_fd_sc_hd__mux2_1
XFILLER_0_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_5_26__f_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_5_26__leaf_clk sky130_fd_sc_hd__clkbuf_16
Xhold2550 data_array.data1\[14\]\[50\] VGND VGND VPWR VPWR net4201 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2561 data_array.data1\[14\]\[32\] VGND VGND VPWR VPWR net4212 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2572 data_array.data1\[3\]\[47\] VGND VGND VPWR VPWR net4223 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2583 data_array.data1\[3\]\[18\] VGND VGND VPWR VPWR net4234 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2594 data_array.data0\[13\]\[1\] VGND VGND VPWR VPWR net4245 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_124_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1860 data_array.data1\[5\]\[60\] VGND VGND VPWR VPWR net3511 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1871 tag_array.tag0\[7\]\[22\] VGND VGND VPWR VPWR net3522 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1882 tag_array.tag1\[6\]\[17\] VGND VGND VPWR VPWR net3533 sky130_fd_sc_hd__dlygate4sd3_1
X_11982_ clknet_leaf_12_clk _00790_ VGND VGND VPWR VPWR data_array.data0\[4\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_91_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1893 tag_array.tag0\[0\]\[15\] VGND VGND VPWR VPWR net3544 sky130_fd_sc_hd__dlygate4sd3_1
X_13721_ clknet_leaf_254_clk _02350_ VGND VGND VPWR VPWR data_array.data1\[1\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_158_3405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10933_ net1008 net4240 net526 VGND VGND VPWR VPWR _02678_ sky130_fd_sc_hd__mux2_1
XFILLER_16_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10864_ net1030 net3529 net524 VGND VGND VPWR VPWR _02609_ sky130_fd_sc_hd__mux2_1
X_13652_ clknet_leaf_85_clk _02281_ VGND VGND VPWR VPWR data_array.data1\[15\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_175_3730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12603_ clknet_leaf_105_clk _01297_ VGND VGND VPWR VPWR tag_array.tag0\[0\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_10795_ net1891 net1051 net508 VGND VGND VPWR VPWR _02540_ sky130_fd_sc_hd__mux2_1
XFILLER_13_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13583_ clknet_leaf_16_clk _02212_ VGND VGND VPWR VPWR data_array.data0\[9\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_171_3638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12534_ clknet_leaf_136_clk _01228_ VGND VGND VPWR VPWR tag_array.tag1\[11\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_171_3649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_928 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12465_ clknet_leaf_254_clk _01159_ VGND VGND VPWR VPWR data_array.data1\[9\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_438 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14204_ clknet_leaf_223_clk _02833_ VGND VGND VPWR VPWR data_array.data0\[2\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
X_11416_ clknet_leaf_210_clk _00226_ VGND VGND VPWR VPWR data_array.data0\[0\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_12396_ clknet_leaf_51_clk _01090_ VGND VGND VPWR VPWR data_array.data0\[14\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_153_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11347_ net906 net4382 net795 VGND VGND VPWR VPWR _03090_ sky130_fd_sc_hd__mux2_1
X_14135_ clknet_leaf_39_clk _02764_ VGND VGND VPWR VPWR data_array.data0\[1\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11278_ net919 net4571 net681 VGND VGND VPWR VPWR _03021_ sky130_fd_sc_hd__mux2_1
X_14066_ clknet_leaf_87_clk _02695_ VGND VGND VPWR VPWR data_array.data1\[6\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
X_13017_ clknet_leaf_260_clk _01711_ VGND VGND VPWR VPWR data_array.data0\[3\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
X_10229_ net889 net4606 net355 VGND VGND VPWR VPWR _01976_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05770_ net20 fsm.tag_out1\[20\] VGND VGND VPWR VPWR _03287_ sky130_fd_sc_hd__or2_1
X_13919_ clknet_leaf_203_clk _02548_ VGND VGND VPWR VPWR data_array.data1\[4\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_18_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07440_ _04680_ _04681_ VGND VGND VPWR VPWR _00059_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07371_ data_array.data0\[4\]\[57\] net1347 net1253 data_array.data0\[7\]\[57\] _04618_
+ VGND VGND VPWR VPWR _04619_ sky130_fd_sc_hd__a221o_1
X_09110_ net1100 net4110 net567 VGND VGND VPWR VPWR _00864_ sky130_fd_sc_hd__mux2_1
X_06322_ tag_array.tag0\[4\]\[12\] net1407 net1313 tag_array.tag0\[7\]\[12\] _03664_
+ VGND VGND VPWR VPWR _03665_ sky130_fd_sc_hd__a221o_1
XFILLER_176_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09041_ net2269 net860 net425 VGND VGND VPWR VPWR _00796_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_96_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06253_ tag_array.tag0\[13\]\[6\] net1597 net1501 tag_array.tag0\[14\]\[6\] VGND
+ VGND VPWR VPWR _03602_ sky130_fd_sc_hd__a22o_1
XFILLER_129_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold401 data_array.data0\[8\]\[63\] VGND VGND VPWR VPWR net2052 sky130_fd_sc_hd__dlygate4sd3_1
X_06184_ net1199 _03533_ _03537_ net1625 VGND VGND VPWR VPWR _03540_ sky130_fd_sc_hd__a22o_1
XFILLER_116_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold412 data_array.data0\[4\]\[55\] VGND VGND VPWR VPWR net2063 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold423 data_array.data1\[1\]\[41\] VGND VGND VPWR VPWR net2074 sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 data_array.data0\[2\]\[53\] VGND VGND VPWR VPWR net2085 sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 data_array.data1\[0\]\[0\] VGND VGND VPWR VPWR net2096 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold456 data_array.data0\[2\]\[51\] VGND VGND VPWR VPWR net2107 sky130_fd_sc_hd__dlygate4sd3_1
Xhold467 data_array.data0\[8\]\[47\] VGND VGND VPWR VPWR net2118 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold478 data_array.data0\[4\]\[30\] VGND VGND VPWR VPWR net2129 sky130_fd_sc_hd__dlygate4sd3_1
Xhold489 data_array.data1\[1\]\[63\] VGND VGND VPWR VPWR net2140 sky130_fd_sc_hd__dlygate4sd3_1
X_09943_ net1058 net3041 net372 VGND VGND VPWR VPWR _01692_ sky130_fd_sc_hd__mux2_1
Xfanout903 _05524_ VGND VGND VPWR VPWR net903 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout914 net915 VGND VGND VPWR VPWR net914 sky130_fd_sc_hd__clkbuf_2
Xfanout925 _05512_ VGND VGND VPWR VPWR net925 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_70_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout936 net939 VGND VGND VPWR VPWR net936 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_70_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout947 _05502_ VGND VGND VPWR VPWR net947 sky130_fd_sc_hd__clkbuf_2
X_09874_ net973 net2847 net378 VGND VGND VPWR VPWR _01624_ sky130_fd_sc_hd__mux2_1
XFILLER_98_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout958 net959 VGND VGND VPWR VPWR net958 sky130_fd_sc_hd__clkbuf_2
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout969 _05490_ VGND VGND VPWR VPWR net969 sky130_fd_sc_hd__buf_1
Xhold1101 tag_array.tag0\[1\]\[13\] VGND VGND VPWR VPWR net2752 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1112 data_array.data0\[2\]\[11\] VGND VGND VPWR VPWR net2763 sky130_fd_sc_hd__dlygate4sd3_1
X_08825_ net2029 net945 net443 VGND VGND VPWR VPWR _00583_ sky130_fd_sc_hd__mux2_1
Xhold1123 tag_array.tag0\[2\]\[18\] VGND VGND VPWR VPWR net2774 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1134 tag_array.tag0\[5\]\[22\] VGND VGND VPWR VPWR net2785 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1145 tag_array.tag1\[12\]\[12\] VGND VGND VPWR VPWR net2796 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1156 tag_array.tag1\[13\]\[24\] VGND VGND VPWR VPWR net2807 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1167 data_array.data1\[15\]\[56\] VGND VGND VPWR VPWR net2818 sky130_fd_sc_hd__dlygate4sd3_1
X_08756_ net701 net3388 net464 VGND VGND VPWR VPWR _00515_ sky130_fd_sc_hd__mux2_1
Xhold1178 tag_array.tag1\[11\]\[4\] VGND VGND VPWR VPWR net2829 sky130_fd_sc_hd__dlygate4sd3_1
X_05968_ net138 net1151 _03438_ _03439_ VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__a22o_1
XFILLER_73_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1189 data_array.data0\[9\]\[6\] VGND VGND VPWR VPWR net2840 sky130_fd_sc_hd__dlygate4sd3_1
X_07707_ data_array.data1\[5\]\[24\] net1577 net1481 data_array.data1\[6\]\[24\] VGND
+ VGND VPWR VPWR _04924_ sky130_fd_sc_hd__a22o_1
X_08687_ net2156 net775 net481 VGND VGND VPWR VPWR _00446_ sky130_fd_sc_hd__mux2_1
X_05899_ net113 net1151 _03392_ _03393_ VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_68_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07638_ _04860_ _04861_ VGND VGND VPWR VPWR _00072_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_68_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07569_ data_array.data1\[4\]\[11\] net1384 net1290 data_array.data1\[7\]\[11\] _04798_
+ VGND VGND VPWR VPWR _04799_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_153_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_153_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09308_ net747 net2658 net553 VGND VGND VPWR VPWR _01062_ sky130_fd_sc_hd__mux2_1
X_10580_ net887 net2818 net455 VGND VGND VPWR VPWR _02325_ sky130_fd_sc_hd__mux2_1
XFILLER_10_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09239_ net722 net3022 net646 VGND VGND VPWR VPWR _00993_ sky130_fd_sc_hd__mux2_1
XFILLER_182_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12250_ clknet_leaf_132_clk _01008_ VGND VGND VPWR VPWR tag_array.tag1\[14\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_11201_ net969 net3774 net648 VGND VGND VPWR VPWR _02944_ sky130_fd_sc_hd__mux2_1
XFILLER_181_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12181_ clknet_leaf_145_clk _00989_ VGND VGND VPWR VPWR tag_array.tag0\[14\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11132_ net991 net2892 net549 VGND VGND VPWR VPWR _02875_ sky130_fd_sc_hd__mux2_1
XFILLER_79_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold990 data_array.data0\[12\]\[26\] VGND VGND VPWR VPWR net2641 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_62_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11063_ net1951 net1009 net328 VGND VGND VPWR VPWR _02806_ sky130_fd_sc_hd__mux2_1
X_10014_ net1030 net3031 net564 VGND VGND VPWR VPWR _01763_ sky130_fd_sc_hd__mux2_1
XFILLER_62_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_129_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2380 data_array.data1\[14\]\[19\] VGND VGND VPWR VPWR net4031 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2391 data_array.data1\[6\]\[7\] VGND VGND VPWR VPWR net4042 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_4_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1690 data_array.data0\[6\]\[38\] VGND VGND VPWR VPWR net3341 sky130_fd_sc_hd__dlygate4sd3_1
X_11965_ clknet_leaf_235_clk _00773_ VGND VGND VPWR VPWR data_array.data0\[4\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13704_ clknet_leaf_227_clk _02333_ VGND VGND VPWR VPWR data_array.data1\[1\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_45_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10916_ net1078 net3209 net531 VGND VGND VPWR VPWR _02661_ sky130_fd_sc_hd__mux2_1
XFILLER_44_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11896_ clknet_leaf_11_clk _00704_ VGND VGND VPWR VPWR data_array.data0\[5\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
X_13635_ clknet_leaf_114_clk _02264_ VGND VGND VPWR VPWR data_array.data0\[9\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
X_10847_ net1098 net3490 net519 VGND VGND VPWR VPWR _02592_ sky130_fd_sc_hd__mux2_1
XFILLER_13_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13566_ clknet_leaf_193_clk _02195_ VGND VGND VPWR VPWR data_array.data1\[0\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
X_10778_ net862 net2969 net500 VGND VGND VPWR VPWR _02523_ sky130_fd_sc_hd__mux2_1
X_12517_ clknet_leaf_178_clk _01211_ VGND VGND VPWR VPWR lru_array.lru_mem\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_74_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13497_ clknet_leaf_35_clk _02126_ VGND VGND VPWR VPWR tag_array.dirty1\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_172_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12448_ clknet_leaf_174_clk _01142_ VGND VGND VPWR VPWR data_array.data1\[9\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12379_ clknet_leaf_201_clk _00057_ VGND VGND VPWR VPWR data_array.rdata0\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_181_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14118_ clknet_leaf_71_clk _02747_ VGND VGND VPWR VPWR data_array.data0\[1\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06940_ data_array.data0\[12\]\[18\] net1343 net1249 data_array.data0\[15\]\[18\]
+ _04226_ VGND VGND VPWR VPWR _04227_ sky130_fd_sc_hd__a221o_1
X_14049_ clknet_leaf_269_clk _02678_ VGND VGND VPWR VPWR data_array.data1\[6\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_68_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06871_ data_array.data0\[1\]\[12\] net1579 net1483 data_array.data0\[2\]\[12\] VGND
+ VGND VPWR VPWR _04164_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_2_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_230_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_230_clk
+ sky130_fd_sc_hd__clkbuf_8
X_08610_ net782 net3866 net518 VGND VGND VPWR VPWR _00369_ sky130_fd_sc_hd__mux2_1
X_05822_ _03139_ fsm.tag_out1\[11\] _03243_ VGND VGND VPWR VPWR _03339_ sky130_fd_sc_hd__o21ai_1
X_09590_ net988 net4580 net399 VGND VGND VPWR VPWR _01342_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_89_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_84_Right_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05753_ net30 fsm.tag_out1\[0\] VGND VGND VPWR VPWR _03270_ sky130_fd_sc_hd__and2b_1
X_08541_ net792 net3436 net585 VGND VGND VPWR VPWR _00309_ sky130_fd_sc_hd__mux2_1
XFILLER_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08472_ _05550_ net815 VGND VGND VPWR VPWR _05551_ sky130_fd_sc_hd__nand2b_4
X_05684_ net8 fsm.tag_out0\[9\] VGND VGND VPWR VPWR _03201_ sky130_fd_sc_hd__and2b_1
XFILLER_165_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07423_ data_array.data0\[13\]\[62\] net1602 net1506 data_array.data0\[14\]\[62\]
+ VGND VGND VPWR VPWR _04666_ sky130_fd_sc_hd__a22o_1
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07354_ data_array.data0\[12\]\[56\] net1342 net1248 data_array.data0\[15\]\[56\]
+ _04602_ VGND VGND VPWR VPWR _04603_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_63_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_114_Left_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06305_ net1207 _03643_ _03647_ net1633 VGND VGND VPWR VPWR _03650_ sky130_fd_sc_hd__a22o_1
XFILLER_149_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07285_ net1226 _04535_ _04539_ net1178 VGND VGND VPWR VPWR _04541_ sky130_fd_sc_hd__a22o_1
XFILLER_108_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09024_ net2402 net928 net419 VGND VGND VPWR VPWR _00779_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_93_Right_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06236_ tag_array.tag0\[12\]\[4\] net1373 net1279 tag_array.tag0\[15\]\[4\] _03586_
+ VGND VGND VPWR VPWR _03587_ sky130_fd_sc_hd__a221o_1
Xhold220 data_array.data1\[4\]\[1\] VGND VGND VPWR VPWR net1871 sky130_fd_sc_hd__dlygate4sd3_1
X_06167_ tag_array.valid0\[13\] net1597 net1501 tag_array.valid0\[14\] VGND VGND VPWR
+ VPWR _03524_ sky130_fd_sc_hd__a22o_1
XFILLER_145_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold231 data_array.data0\[4\]\[17\] VGND VGND VPWR VPWR net1882 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold242 data_array.data0\[4\]\[46\] VGND VGND VPWR VPWR net1893 sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 data_array.data1\[0\]\[55\] VGND VGND VPWR VPWR net1904 sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 data_array.data0\[1\]\[8\] VGND VGND VPWR VPWR net1915 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06098_ data_array.rdata0\[13\] net1136 net1117 data_array.rdata1\[13\] VGND VGND
+ VPWR VPWR net267 sky130_fd_sc_hd__a22o_1
Xhold275 data_array.data0\[1\]\[56\] VGND VGND VPWR VPWR net1926 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout700 net701 VGND VGND VPWR VPWR net700 sky130_fd_sc_hd__clkbuf_2
XFILLER_104_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold286 data_array.data1\[8\]\[49\] VGND VGND VPWR VPWR net1937 sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 data_array.data1\[8\]\[30\] VGND VGND VPWR VPWR net1948 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout711 _05405_ VGND VGND VPWR VPWR net711 sky130_fd_sc_hd__dlymetal6s2s_1
X_09926_ net704 net3106 net604 VGND VGND VPWR VPWR _01676_ sky130_fd_sc_hd__mux2_1
Xfanout722 net723 VGND VGND VPWR VPWR net722 sky130_fd_sc_hd__clkbuf_2
XFILLER_132_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout733 _05395_ VGND VGND VPWR VPWR net733 sky130_fd_sc_hd__buf_1
Xfanout744 net745 VGND VGND VPWR VPWR net744 sky130_fd_sc_hd__clkbuf_2
Xfanout755 _05383_ VGND VGND VPWR VPWR net755 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout766 net767 VGND VGND VPWR VPWR net766 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_146_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09857_ net1042 net4047 net380 VGND VGND VPWR VPWR _01607_ sky130_fd_sc_hd__mux2_1
Xfanout777 _05373_ VGND VGND VPWR VPWR net777 sky130_fd_sc_hd__buf_1
Xfanout788 net790 VGND VGND VPWR VPWR net788 sky130_fd_sc_hd__buf_1
Xfanout799 net806 VGND VGND VPWR VPWR net799 sky130_fd_sc_hd__clkbuf_8
XFILLER_85_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_221_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_221_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_85_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08808_ net2240 net1012 net446 VGND VGND VPWR VPWR _00566_ sky130_fd_sc_hd__mux2_1
XFILLER_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_107_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09788_ net1059 net3417 net388 VGND VGND VPWR VPWR _01539_ sky130_fd_sc_hd__mux2_1
XFILLER_27_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08739_ net766 net3040 net458 VGND VGND VPWR VPWR _00498_ sky130_fd_sc_hd__mux2_1
XFILLER_121_20 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11750_ clknet_leaf_224_clk _00558_ VGND VGND VPWR VPWR data_array.data0\[8\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_92_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10701_ net2153 net914 net484 VGND VGND VPWR VPWR _02446_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_120_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ clknet_leaf_197_clk _00489_ VGND VGND VPWR VPWR tag_array.tag1\[1\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_13420_ clknet_leaf_122_clk _02050_ VGND VGND VPWR VPWR data_array.data1\[8\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
X_10632_ net1748 net934 net473 VGND VGND VPWR VPWR _02377_ sky130_fd_sc_hd__mux2_1
X_13351_ clknet_leaf_115_clk _01981_ VGND VGND VPWR VPWR data_array.data0\[10\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
X_10563_ net953 net4273 net456 VGND VGND VPWR VPWR _02308_ sky130_fd_sc_hd__mux2_1
XFILLER_127_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12302_ clknet_leaf_127_clk _01060_ VGND VGND VPWR VPWR tag_array.tag1\[12\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_127_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10494_ net970 net2364 net345 VGND VGND VPWR VPWR _02239_ sky130_fd_sc_hd__mux2_1
X_13282_ clknet_leaf_13_clk _01912_ VGND VGND VPWR VPWR data_array.data0\[11\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_20_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12233_ clknet_leaf_151_clk _00162_ VGND VGND VPWR VPWR fsm.tag_out1\[15\] sky130_fd_sc_hd__dfxtp_1
X_12164_ clknet_leaf_155_clk _00972_ VGND VGND VPWR VPWR tag_array.tag0\[13\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_166_3548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11115_ net1056 net2619 net545 VGND VGND VPWR VPWR _02858_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12095_ clknet_leaf_258_clk _00903_ VGND VGND VPWR VPWR data_array.data1\[14\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_111_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_183_3873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_3884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11046_ net2574 net1076 net329 VGND VGND VPWR VPWR _02789_ sky130_fd_sc_hd__mux2_1
XFILLER_103_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_212_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_212_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_162_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12997_ clknet_leaf_94_clk _01691_ VGND VGND VPWR VPWR data_array.data0\[3\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_73_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11948_ clknet_leaf_8_clk _00756_ VGND VGND VPWR VPWR data_array.data0\[4\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_11879_ clknet_leaf_249_clk _00687_ VGND VGND VPWR VPWR data_array.data0\[5\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13618_ clknet_leaf_46_clk _02247_ VGND VGND VPWR VPWR data_array.data0\[9\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_38_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13549_ clknet_leaf_261_clk _02178_ VGND VGND VPWR VPWR data_array.data1\[0\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_146_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07070_ data_array.data0\[4\]\[30\] net1392 net1298 data_array.data0\[7\]\[30\] _04344_
+ VGND VGND VPWR VPWR _04345_ sky130_fd_sc_hd__a221o_1
XFILLER_134_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06021_ data_array.rdata1\[63\] net831 net839 VGND VGND VPWR VPWR _03475_ sky130_fd_sc_hd__a21o_1
Xoutput303 net303 VGND VGND VPWR VPWR mem_wdata[46] sky130_fd_sc_hd__buf_2
Xoutput314 net314 VGND VGND VPWR VPWR mem_wdata[56] sky130_fd_sc_hd__buf_2
XFILLER_127_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput325 net325 VGND VGND VPWR VPWR mem_wdata[8] sky130_fd_sc_hd__buf_2
XFILLER_59_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07972_ data_array.data1\[4\]\[48\] net1393 net1299 data_array.data1\[7\]\[48\] _05164_
+ VGND VGND VPWR VPWR _05165_ sky130_fd_sc_hd__a221o_1
XFILLER_101_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09711_ net744 net2584 net609 VGND VGND VPWR VPWR _01463_ sky130_fd_sc_hd__mux2_1
X_06923_ _04210_ _04211_ VGND VGND VPWR VPWR _00007_ sky130_fd_sc_hd__or2_1
XFILLER_67_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_203_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_203_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_67_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09642_ net719 net2638 net615 VGND VGND VPWR VPWR _01394_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06854_ data_array.data0\[0\]\[10\] net1411 net1317 data_array.data0\[3\]\[10\] _04148_
+ VGND VGND VPWR VPWR _04149_ sky130_fd_sc_hd__a221o_1
XFILLER_83_745 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05805_ fsm.tag_out0\[23\] net24 VGND VGND VPWR VPWR _03322_ sky130_fd_sc_hd__and2b_1
X_06785_ data_array.data0\[13\]\[4\] net1582 net1486 data_array.data0\[14\]\[4\] VGND
+ VGND VPWR VPWR _04086_ sky130_fd_sc_hd__a22o_1
X_09573_ net1059 net3963 net396 VGND VGND VPWR VPWR _01325_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_141_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08524_ _03509_ _03519_ VGND VGND VPWR VPWR _05587_ sky130_fd_sc_hd__nor2_1
X_05736_ _03249_ _03250_ _03251_ _03252_ VGND VGND VPWR VPWR _03253_ sky130_fd_sc_hd__or4_1
XFILLER_36_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08455_ net1129 _05539_ VGND VGND VPWR VPWR _05540_ sky130_fd_sc_hd__and2_1
X_05667_ fsm.tag_out0\[16\] net16 VGND VGND VPWR VPWR _03184_ sky130_fd_sc_hd__and2b_1
XFILLER_24_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_82_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_122_Left_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07406_ net1183 _04645_ _04649_ net1231 VGND VGND VPWR VPWR _04651_ sky130_fd_sc_hd__a22o_1
XFILLER_149_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08386_ net1125 _05493_ VGND VGND VPWR VPWR _05494_ sky130_fd_sc_hd__and2_1
XFILLER_91_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07337_ data_array.data0\[5\]\[54\] net1547 net1451 data_array.data0\[6\]\[54\] VGND
+ VGND VPWR VPWR _04588_ sky130_fd_sc_hd__a22o_1
XFILLER_183_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_883 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07268_ data_array.data0\[4\]\[48\] net1387 net1293 data_array.data0\[7\]\[48\] _04524_
+ VGND VGND VPWR VPWR _04525_ sky130_fd_sc_hd__a221o_1
XFILLER_137_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09007_ net2452 net996 net419 VGND VGND VPWR VPWR _00762_ sky130_fd_sc_hd__mux2_1
X_06219_ _03570_ _03571_ VGND VGND VPWR VPWR _00148_ sky130_fd_sc_hd__or2_1
XFILLER_124_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07199_ data_array.data0\[9\]\[42\] net1579 net1483 data_array.data0\[10\]\[42\]
+ VGND VGND VPWR VPWR _04462_ sky130_fd_sc_hd__a22o_1
XFILLER_183_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_148_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_131_Left_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1506 net1507 VGND VGND VPWR VPWR net1506 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1517 net1518 VGND VGND VPWR VPWR net1517 sky130_fd_sc_hd__clkbuf_4
Xfanout1528 net1529 VGND VGND VPWR VPWR net1528 sky130_fd_sc_hd__clkbuf_4
Xfanout530 _05598_ VGND VGND VPWR VPWR net530 sky130_fd_sc_hd__clkbuf_8
Xfanout541 net547 VGND VGND VPWR VPWR net541 sky130_fd_sc_hd__buf_4
Xfanout1539 net1543 VGND VGND VPWR VPWR net1539 sky130_fd_sc_hd__clkbuf_2
Xfanout552 net553 VGND VGND VPWR VPWR net552 sky130_fd_sc_hd__clkbuf_4
X_09909_ net770 net3919 net603 VGND VGND VPWR VPWR _01659_ sky130_fd_sc_hd__mux2_1
Xfanout563 _05593_ VGND VGND VPWR VPWR net563 sky130_fd_sc_hd__buf_4
Xfanout574 net575 VGND VGND VPWR VPWR net574 sky130_fd_sc_hd__buf_4
XFILLER_19_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout585 net590 VGND VGND VPWR VPWR net585 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_161_3456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12920_ clknet_leaf_97_clk _01614_ VGND VGND VPWR VPWR data_array.data0\[13\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout596 net598 VGND VGND VPWR VPWR net596 sky130_fd_sc_hd__buf_4
XFILLER_58_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12851_ clknet_leaf_59_clk _01545_ VGND VGND VPWR VPWR data_array.data0\[12\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_122_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11802_ clknet_leaf_72_clk _00610_ VGND VGND VPWR VPWR data_array.data0\[7\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12782_ clknet_leaf_96_clk _01476_ VGND VGND VPWR VPWR tag_array.tag1\[10\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_140_Left_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11733_ clknet_leaf_185_clk _00541_ VGND VGND VPWR VPWR tag_array.tag0\[9\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_148_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ clknet_leaf_117_clk _03075_ VGND VGND VPWR VPWR data_array.data1\[7\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_175_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11664_ clknet_leaf_135_clk _00472_ VGND VGND VPWR VPWR tag_array.tag1\[1\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_13403_ clknet_leaf_193_clk _02033_ VGND VGND VPWR VPWR data_array.data1\[8\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_10615_ net2225 net1000 net468 VGND VGND VPWR VPWR _02360_ sky130_fd_sc_hd__mux2_1
X_14383_ clknet_leaf_77_clk _03006_ VGND VGND VPWR VPWR data_array.data1\[10\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11595_ clknet_leaf_33_clk _00403_ VGND VGND VPWR VPWR tag_array.tag1\[4\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_167_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13334_ clknet_leaf_46_clk _01964_ VGND VGND VPWR VPWR data_array.data0\[10\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
X_10546_ net1023 net3617 net455 VGND VGND VPWR VPWR _02291_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_137_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13265_ clknet_leaf_88_clk _01895_ VGND VGND VPWR VPWR data_array.data0\[11\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
X_10477_ net1037 net3208 net348 VGND VGND VPWR VPWR _02222_ sky130_fd_sc_hd__mux2_1
X_12216_ clknet_leaf_146_clk _00146_ VGND VGND VPWR VPWR fsm.tag_out0\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_155_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13196_ clknet_leaf_77_clk _00090_ VGND VGND VPWR VPWR data_array.rdata1\[33\] sky130_fd_sc_hd__dfxtp_1
X_12147_ clknet_leaf_178_clk _00955_ VGND VGND VPWR VPWR tag_array.tag0\[13\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_97_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12078_ clknet_leaf_93_clk _00886_ VGND VGND VPWR VPWR data_array.data1\[14\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_77_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11029_ net1926 net884 net337 VGND VGND VPWR VPWR _02773_ sky130_fd_sc_hd__mux2_1
XFILLER_110_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06570_ net1184 _03885_ _03889_ net1232 VGND VGND VPWR VPWR _03891_ sky130_fd_sc_hd__a22o_1
XFILLER_45_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08240_ fsm.tag_out1\[15\] net818 net810 fsm.tag_out0\[15\] _05394_ VGND VGND VPWR
+ VPWR _05395_ sky130_fd_sc_hd__a221o_2
XFILLER_60_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_15 _03133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_26 _05405_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_37 net393 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_48 net666 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08171_ lru_array.lru_mem\[9\] net1564 net1468 lru_array.lru_mem\[10\] VGND VGND
+ VPWR VPWR _05346_ sky130_fd_sc_hd__a22o_1
XANTENNA_59 net1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07122_ data_array.data0\[13\]\[35\] net1537 net1441 data_array.data0\[14\]\[35\]
+ VGND VGND VPWR VPWR _04392_ sky130_fd_sc_hd__a22o_1
XFILLER_146_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07053_ net1619 _04323_ _04327_ net1193 VGND VGND VPWR VPWR _04330_ sky130_fd_sc_hd__a22o_1
XFILLER_134_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06004_ net151 net1152 _03462_ _03463_ VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__a22o_1
XFILLER_114_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput166 net166 VGND VGND VPWR VPWR cpu_rdata[10] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_58_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput177 net177 VGND VGND VPWR VPWR cpu_rdata[20] sky130_fd_sc_hd__buf_2
Xoutput188 net188 VGND VGND VPWR VPWR cpu_rdata[30] sky130_fd_sc_hd__buf_6
XFILLER_130_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2902 data_array.data1\[6\]\[54\] VGND VGND VPWR VPWR net4553 sky130_fd_sc_hd__dlygate4sd3_1
Xoutput199 net199 VGND VGND VPWR VPWR cpu_rdata[40] sky130_fd_sc_hd__buf_2
Xclkbuf_5_7__f_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_5_7__leaf_clk sky130_fd_sc_hd__clkbuf_16
Xhold2913 data_array.data0\[6\]\[31\] VGND VGND VPWR VPWR net4564 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_141_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2924 data_array.data1\[10\]\[33\] VGND VGND VPWR VPWR net4575 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2935 data_array.data1\[11\]\[53\] VGND VGND VPWR VPWR net4586 sky130_fd_sc_hd__dlygate4sd3_1
X_07955_ net1614 _05143_ _05147_ net1189 VGND VGND VPWR VPWR _05150_ sky130_fd_sc_hd__a22o_1
XFILLER_130_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2946 tag_array.tag1\[7\]\[9\] VGND VGND VPWR VPWR net4597 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2957 tag_array.tag1\[14\]\[0\] VGND VGND VPWR VPWR net4608 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_143_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2968 data_array.data0\[13\]\[28\] VGND VGND VPWR VPWR net4619 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_101_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06906_ data_array.data0\[13\]\[15\] net1580 net1484 data_array.data0\[14\]\[15\]
+ VGND VGND VPWR VPWR _04196_ sky130_fd_sc_hd__a22o_1
X_07886_ data_array.data1\[8\]\[40\] net1415 net1321 data_array.data1\[11\]\[40\]
+ _05086_ VGND VGND VPWR VPWR _05087_ sky130_fd_sc_hd__a221o_1
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09625_ net789 net2771 net615 VGND VGND VPWR VPWR _01377_ sky130_fd_sc_hd__mux2_1
X_06837_ data_array.data0\[8\]\[9\] net1389 net1295 data_array.data0\[11\]\[9\] _04132_
+ VGND VGND VPWR VPWR _04133_ sky130_fd_sc_hd__a221o_1
X_09556_ net705 net2349 net620 VGND VGND VPWR VPWR _01309_ sky130_fd_sc_hd__mux2_1
X_06768_ net1166 _04065_ _04069_ net1215 VGND VGND VPWR VPWR _04071_ sky130_fd_sc_hd__a22o_1
X_08507_ _03511_ _03527_ net822 VGND VGND VPWR VPWR _05575_ sky130_fd_sc_hd__or3_1
XFILLER_169_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05719_ _03217_ _03226_ _03231_ _03235_ VGND VGND VPWR VPWR _03236_ sky130_fd_sc_hd__nor4_1
XFILLER_70_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09487_ net781 net3061 net624 VGND VGND VPWR VPWR _01240_ sky130_fd_sc_hd__mux2_1
X_06699_ tag_array.tag1\[1\]\[21\] net1592 net1496 tag_array.tag1\[2\]\[21\] VGND
+ VGND VPWR VPWR _04008_ sky130_fd_sc_hd__a22o_1
XFILLER_178_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08438_ net3004 net895 net688 VGND VGND VPWR VPWR _00275_ sky130_fd_sc_hd__mux2_1
XFILLER_169_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08369_ net1820 net986 net692 VGND VGND VPWR VPWR _00252_ sky130_fd_sc_hd__mux2_1
XFILLER_149_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10400_ net2036 net1055 net667 VGND VGND VPWR VPWR _02146_ sky130_fd_sc_hd__mux2_1
XFILLER_183_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11380_ net164 VGND VGND VPWR VPWR _00190_ sky130_fd_sc_hd__inv_2
XFILLER_164_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10331_ net776 net3808 net591 VGND VGND VPWR VPWR _02078_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_115_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13050_ clknet_leaf_264_clk _01744_ VGND VGND VPWR VPWR data_array.data1\[13\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_10262_ net694 net2308 net595 VGND VGND VPWR VPWR _02009_ sky130_fd_sc_hd__mux2_1
XFILLER_124_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12001_ clknet_leaf_45_clk _00809_ VGND VGND VPWR VPWR data_array.data0\[6\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_79_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10193_ net1032 net2882 net359 VGND VGND VPWR VPWR _01940_ sky130_fd_sc_hd__mux2_1
XFILLER_120_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1303 net1304 VGND VGND VPWR VPWR net1303 sky130_fd_sc_hd__clkbuf_4
Xfanout1314 net1328 VGND VGND VPWR VPWR net1314 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_180_3810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1325 net1326 VGND VGND VPWR VPWR net1325 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_180_3821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1336 net1339 VGND VGND VPWR VPWR net1336 sky130_fd_sc_hd__clkbuf_4
Xfanout1347 net1348 VGND VGND VPWR VPWR net1347 sky130_fd_sc_hd__clkbuf_4
XFILLER_47_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1358 net1364 VGND VGND VPWR VPWR net1358 sky130_fd_sc_hd__clkbuf_2
Xfanout360 net361 VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__clkbuf_8
Xfanout371 net374 VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__buf_4
Xfanout1369 net1370 VGND VGND VPWR VPWR net1369 sky130_fd_sc_hd__clkbuf_4
Xfanout382 net384 VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__clkbuf_8
Xfanout393 _03125_ VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__clkbuf_8
X_13952_ clknet_leaf_21_clk _02581_ VGND VGND VPWR VPWR data_array.data1\[4\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12903_ clknet_leaf_104_clk _01597_ VGND VGND VPWR VPWR data_array.data0\[13\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_13883_ clknet_leaf_4_clk _02512_ VGND VGND VPWR VPWR data_array.data1\[3\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12834_ clknet_leaf_248_clk _01528_ VGND VGND VPWR VPWR data_array.data0\[12\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_178_3772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_3783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ clknet_leaf_144_clk _01459_ VGND VGND VPWR VPWR tag_array.tag0\[6\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_11716_ clknet_leaf_143_clk _00524_ VGND VGND VPWR VPWR tag_array.tag0\[9\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12696_ clknet_leaf_173_clk _01390_ VGND VGND VPWR VPWR tag_array.tag0\[8\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14435_ clknet_leaf_66_clk _03058_ VGND VGND VPWR VPWR data_array.data1\[7\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_11647_ clknet_leaf_133_clk _00455_ VGND VGND VPWR VPWR tag_array.tag1\[2\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput13 cpu_addr[20] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_2
XFILLER_174_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput24 cpu_addr[30] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_2
Xinput35 cpu_wdata[10] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_1
X_14366_ clknet_leaf_213_clk _02989_ VGND VGND VPWR VPWR data_array.data1\[10\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput46 cpu_wdata[20] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_1
X_11578_ clknet_leaf_98_clk _00386_ VGND VGND VPWR VPWR tag_array.tag1\[5\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput57 cpu_wdata[30] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_1
Xinput68 cpu_wdata[40] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_1
XFILLER_171_812 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold808 data_array.data0\[12\]\[19\] VGND VGND VPWR VPWR net2459 sky130_fd_sc_hd__dlygate4sd3_1
X_13317_ clknet_leaf_245_clk _01947_ VGND VGND VPWR VPWR data_array.data0\[10\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_10529_ net1091 net3876 net457 VGND VGND VPWR VPWR _02274_ sky130_fd_sc_hd__mux2_1
Xinput79 cpu_wdata[50] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_1
Xhold819 data_array.data0\[7\]\[26\] VGND VGND VPWR VPWR net2470 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_172_Right_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14297_ clknet_leaf_254_clk _02926_ VGND VGND VPWR VPWR data_array.data1\[11\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_109_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13248_ clknet_leaf_228_clk _01878_ VGND VGND VPWR VPWR data_array.data0\[11\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_170_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13179_ clknet_leaf_212_clk _00071_ VGND VGND VPWR VPWR data_array.rdata1\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_124_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2209 data_array.data1\[15\]\[18\] VGND VGND VPWR VPWR net3860 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_36_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1508 data_array.data0\[2\]\[14\] VGND VGND VPWR VPWR net3159 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1519 data_array.data1\[14\]\[28\] VGND VGND VPWR VPWR net3170 sky130_fd_sc_hd__dlygate4sd3_1
X_07740_ data_array.data1\[1\]\[27\] net1528 net1432 data_array.data1\[2\]\[27\] VGND
+ VGND VPWR VPWR _04954_ sky130_fd_sc_hd__a22o_1
X_07671_ _04890_ _04891_ VGND VGND VPWR VPWR _00076_ sky130_fd_sc_hd__or2_1
XFILLER_37_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09410_ net1024 net3575 net582 VGND VGND VPWR VPWR _01163_ sky130_fd_sc_hd__mux2_1
X_06622_ tag_array.tag1\[5\]\[14\] net1558 net1462 tag_array.tag1\[6\]\[14\] VGND
+ VGND VPWR VPWR _03938_ sky130_fd_sc_hd__a22o_1
X_06553_ tag_array.tag1\[4\]\[8\] net1417 net1323 tag_array.tag1\[7\]\[8\] _03874_
+ VGND VGND VPWR VPWR _03875_ sky130_fd_sc_hd__a221o_1
X_09341_ net1036 net4199 net403 VGND VGND VPWR VPWR _01094_ sky130_fd_sc_hd__mux2_1
XFILLER_179_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06484_ tag_array.tag1\[9\]\[2\] net1575 net1479 tag_array.tag1\[10\]\[2\] VGND VGND
+ VPWR VPWR _03812_ sky130_fd_sc_hd__a22o_1
X_09272_ net792 net4235 net561 VGND VGND VPWR VPWR _01026_ sky130_fd_sc_hd__mux2_1
XFILLER_179_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08223_ net756 net4597 net804 VGND VGND VPWR VPWR _00205_ sky130_fd_sc_hd__mux2_1
XFILLER_147_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08154_ net1217 _05325_ _05329_ net1169 VGND VGND VPWR VPWR _05331_ sky130_fd_sc_hd__a22o_1
XFILLER_146_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07105_ data_array.data0\[8\]\[33\] net1396 net1302 data_array.data0\[11\]\[33\]
+ _04376_ VGND VGND VPWR VPWR _04377_ sky130_fd_sc_hd__a221o_1
X_08085_ data_array.data1\[1\]\[58\] net1550 net1454 data_array.data1\[2\]\[58\] VGND
+ VGND VPWR VPWR _05268_ sky130_fd_sc_hd__a22o_1
XFILLER_106_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload240 clknet_leaf_137_clk VGND VGND VPWR VPWR clkload240/Y sky130_fd_sc_hd__inv_6
X_07036_ data_array.data0\[1\]\[27\] net1538 net1442 data_array.data0\[2\]\[27\] VGND
+ VGND VPWR VPWR _04314_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_77_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_889 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2710 data_array.data0\[15\]\[17\] VGND VGND VPWR VPWR net4361 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_73_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2721 data_array.data0\[9\]\[23\] VGND VGND VPWR VPWR net4372 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_110_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2732 tag_array.tag1\[6\]\[19\] VGND VGND VPWR VPWR net4383 sky130_fd_sc_hd__dlygate4sd3_1
X_08987_ net1916 net1076 net418 VGND VGND VPWR VPWR _00742_ sky130_fd_sc_hd__mux2_1
Xhold2743 data_array.data0\[7\]\[51\] VGND VGND VPWR VPWR net4394 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_5_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_5_0_clk sky130_fd_sc_hd__clkbuf_8
Xhold2754 tag_array.tag0\[10\]\[23\] VGND VGND VPWR VPWR net4405 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_180_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2765 data_array.data1\[11\]\[59\] VGND VGND VPWR VPWR net4416 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2776 data_array.data0\[3\]\[54\] VGND VGND VPWR VPWR net4427 sky130_fd_sc_hd__dlygate4sd3_1
X_07938_ data_array.data1\[1\]\[45\] net1540 net1444 data_array.data1\[2\]\[45\] VGND
+ VGND VPWR VPWR _05134_ sky130_fd_sc_hd__a22o_1
Xhold2787 data_array.data1\[5\]\[21\] VGND VGND VPWR VPWR net4438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2798 data_array.data1\[11\]\[16\] VGND VGND VPWR VPWR net4449 sky130_fd_sc_hd__dlygate4sd3_1
X_07869_ _05070_ _05071_ VGND VGND VPWR VPWR _00095_ sky130_fd_sc_hd__or2_1
XFILLER_84_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09608_ net916 net3638 net399 VGND VGND VPWR VPWR _01360_ sky130_fd_sc_hd__mux2_1
XFILLER_73_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10880_ net966 net2576 net523 VGND VGND VPWR VPWR _02625_ sky130_fd_sc_hd__mux2_1
X_09539_ net771 net4071 net619 VGND VGND VPWR VPWR _01292_ sky130_fd_sc_hd__mux2_1
XFILLER_25_973 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12550_ clknet_leaf_143_clk _01244_ VGND VGND VPWR VPWR tag_array.tag0\[11\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_156_3355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11501_ clknet_leaf_95_clk _00309_ VGND VGND VPWR VPWR tag_array.tag1\[9\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_12481_ clknet_leaf_76_clk _01175_ VGND VGND VPWR VPWR data_array.data1\[9\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_173_3680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14220_ clknet_leaf_68_clk _02849_ VGND VGND VPWR VPWR data_array.data1\[12\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_156_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11432_ clknet_leaf_226_clk _00242_ VGND VGND VPWR VPWR data_array.data0\[0\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_134_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14151_ clknet_leaf_224_clk _02780_ VGND VGND VPWR VPWR data_array.data0\[1\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
X_11363_ net1648 net2442 net596 VGND VGND VPWR VPWR _03106_ sky130_fd_sc_hd__mux2_1
XFILLER_125_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13102_ clknet_leaf_5_clk _01796_ VGND VGND VPWR VPWR data_array.data1\[13\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
X_10314_ net3349 net906 net633 VGND VGND VPWR VPWR _02061_ sky130_fd_sc_hd__mux2_1
X_14082_ clknet_leaf_201_clk _02711_ VGND VGND VPWR VPWR data_array.data1\[6\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
X_11294_ net820 net3806 _05559_ VGND VGND VPWR VPWR _03037_ sky130_fd_sc_hd__mux2_1
XFILLER_98_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13033_ clknet_leaf_40_clk _01727_ VGND VGND VPWR VPWR data_array.data0\[3\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
X_10245_ net763 net4179 net596 VGND VGND VPWR VPWR _01992_ sky130_fd_sc_hd__mux2_1
XFILLER_26_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1100 _05424_ VGND VGND VPWR VPWR net1100 sky130_fd_sc_hd__clkbuf_2
XFILLER_65_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1111 _05420_ VGND VGND VPWR VPWR net1111 sky130_fd_sc_hd__clkbuf_1
X_10176_ net1103 net2443 net356 VGND VGND VPWR VPWR _01923_ sky130_fd_sc_hd__mux2_1
Xfanout1122 _03478_ VGND VGND VPWR VPWR net1122 sky130_fd_sc_hd__clkbuf_2
XFILLER_78_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1133 _03479_ VGND VGND VPWR VPWR net1133 sky130_fd_sc_hd__buf_2
Xfanout1144 net1145 VGND VGND VPWR VPWR net1144 sky130_fd_sc_hd__clkbuf_4
Xfanout1155 net1156 VGND VGND VPWR VPWR net1155 sky130_fd_sc_hd__buf_4
Xfanout1166 net1167 VGND VGND VPWR VPWR net1166 sky130_fd_sc_hd__buf_4
XFILLER_120_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1177 net1187 VGND VGND VPWR VPWR net1177 sky130_fd_sc_hd__buf_4
Xfanout1188 net1191 VGND VGND VPWR VPWR net1188 sky130_fd_sc_hd__buf_4
Xfanout1199 net1200 VGND VGND VPWR VPWR net1199 sky130_fd_sc_hd__clkbuf_4
X_13935_ clknet_leaf_240_clk _02564_ VGND VGND VPWR VPWR data_array.data1\[4\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_704 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13866_ clknet_leaf_8_clk _02495_ VGND VGND VPWR VPWR data_array.data1\[3\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
X_12817_ clknet_leaf_105_clk _01511_ VGND VGND VPWR VPWR tag_array.tag1\[0\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_13797_ clknet_leaf_40_clk _02426_ VGND VGND VPWR VPWR data_array.data1\[2\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_12748_ clknet_leaf_157_clk _01442_ VGND VGND VPWR VPWR tag_array.tag0\[5\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_148_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12679_ clknet_leaf_205_clk _01373_ VGND VGND VPWR VPWR data_array.data0\[15\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_13_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14418_ clknet_leaf_252_clk _03041_ VGND VGND VPWR VPWR data_array.data1\[7\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14349_ clknet_leaf_184_clk _00185_ _00194_ VGND VGND VPWR VPWR fsm.state\[5\] sky130_fd_sc_hd__dfrtp_1
Xhold605 data_array.data0\[4\]\[29\] VGND VGND VPWR VPWR net2256 sky130_fd_sc_hd__dlygate4sd3_1
Xhold616 data_array.data0\[1\]\[59\] VGND VGND VPWR VPWR net2267 sky130_fd_sc_hd__dlygate4sd3_1
Xhold627 data_array.data0\[0\]\[57\] VGND VGND VPWR VPWR net2278 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold638 tag_array.tag0\[11\]\[14\] VGND VGND VPWR VPWR net2289 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_94_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold649 tag_array.tag1\[8\]\[3\] VGND VGND VPWR VPWR net2300 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_94_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08910_ net866 net3618 net436 VGND VGND VPWR VPWR _00667_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09890_ net909 net4492 net379 VGND VGND VPWR VPWR _01640_ sky130_fd_sc_hd__mux2_1
XFILLER_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2006 tag_array.tag0\[0\]\[6\] VGND VGND VPWR VPWR net3657 sky130_fd_sc_hd__dlygate4sd3_1
X_08841_ net1945 net881 net445 VGND VGND VPWR VPWR _00599_ sky130_fd_sc_hd__mux2_1
Xhold2017 tag_array.tag0\[1\]\[18\] VGND VGND VPWR VPWR net3668 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2028 data_array.data1\[13\]\[45\] VGND VGND VPWR VPWR net3679 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2039 data_array.data0\[11\]\[9\] VGND VGND VPWR VPWR net3690 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1305 tag_array.tag0\[13\]\[20\] VGND VGND VPWR VPWR net2956 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1316 tag_array.tag0\[8\]\[4\] VGND VGND VPWR VPWR net2967 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1327 data_array.data0\[12\]\[48\] VGND VGND VPWR VPWR net2978 sky130_fd_sc_hd__dlygate4sd3_1
X_08772_ net736 net2783 net450 VGND VGND VPWR VPWR _00531_ sky130_fd_sc_hd__mux2_1
X_05984_ data_array.rdata0\[51\] net846 net1142 VGND VGND VPWR VPWR _03450_ sky130_fd_sc_hd__o21a_1
Xhold1338 data_array.data1\[15\]\[16\] VGND VGND VPWR VPWR net2989 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1349 data_array.data1\[7\]\[60\] VGND VGND VPWR VPWR net3000 sky130_fd_sc_hd__dlygate4sd3_1
X_07723_ data_array.data1\[4\]\[25\] net1329 net1235 data_array.data1\[7\]\[25\] _04938_
+ VGND VGND VPWR VPWR _04939_ sky130_fd_sc_hd__a221o_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07654_ data_array.data1\[9\]\[19\] net1584 net1488 data_array.data1\[10\]\[19\]
+ VGND VGND VPWR VPWR _04876_ sky130_fd_sc_hd__a22o_1
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06605_ tag_array.tag1\[13\]\[13\] net1611 net1515 tag_array.tag1\[14\]\[13\] VGND
+ VGND VPWR VPWR _03922_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07585_ data_array.data1\[12\]\[13\] net1364 net1270 data_array.data1\[15\]\[13\]
+ _04812_ VGND VGND VPWR VPWR _04813_ sky130_fd_sc_hd__a221o_1
XFILLER_40_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09324_ net1105 net4602 net402 VGND VGND VPWR VPWR _01077_ sky130_fd_sc_hd__mux2_1
X_06536_ net1197 _03853_ _03857_ net1623 VGND VGND VPWR VPWR _03860_ sky130_fd_sc_hd__a22o_1
XFILLER_159_28 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09255_ net761 net3348 net577 VGND VGND VPWR VPWR _01009_ sky130_fd_sc_hd__mux2_1
X_06467_ tag_array.tag1\[12\]\[0\] net1386 net1292 tag_array.tag1\[15\]\[0\] _03796_
+ VGND VGND VPWR VPWR _03797_ sky130_fd_sc_hd__a221o_1
X_08206_ net1649 net1160 net3 VGND VGND VPWR VPWR _05372_ sky130_fd_sc_hd__and3_1
X_09186_ net736 net2863 net627 VGND VGND VPWR VPWR _00940_ sky130_fd_sc_hd__mux2_1
X_06398_ tag_array.tag0\[1\]\[19\] net1595 net1499 tag_array.tag0\[2\]\[19\] VGND
+ VGND VPWR VPWR _03734_ sky130_fd_sc_hd__a22o_1
XFILLER_147_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08137_ data_array.data1\[4\]\[63\] net1361 net1267 data_array.data1\[7\]\[63\] _05314_
+ VGND VGND VPWR VPWR _05315_ sky130_fd_sc_hd__a221o_1
XFILLER_111_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08068_ data_array.data1\[13\]\[57\] net1538 net1442 data_array.data1\[14\]\[57\]
+ VGND VGND VPWR VPWR _05252_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_112_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07019_ data_array.data0\[4\]\[25\] net1329 net1235 data_array.data0\[7\]\[25\] _04298_
+ VGND VGND VPWR VPWR _04299_ sky130_fd_sc_hd__a221o_1
XFILLER_108_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10030_ net967 net2575 net563 VGND VGND VPWR VPWR _01779_ sky130_fd_sc_hd__mux2_1
XFILLER_0_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2540 data_array.data1\[7\]\[31\] VGND VGND VPWR VPWR net4191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2551 tag_array.tag0\[0\]\[4\] VGND VGND VPWR VPWR net4202 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2562 tag_array.tag0\[12\]\[23\] VGND VGND VPWR VPWR net4213 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2573 data_array.data1\[14\]\[9\] VGND VGND VPWR VPWR net4224 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2584 tag_array.tag1\[13\]\[0\] VGND VGND VPWR VPWR net4235 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2595 data_array.data0\[10\]\[0\] VGND VGND VPWR VPWR net4246 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1850 data_array.data1\[2\]\[31\] VGND VGND VPWR VPWR net3501 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1861 data_array.data1\[10\]\[58\] VGND VGND VPWR VPWR net3512 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1872 tag_array.tag1\[15\]\[13\] VGND VGND VPWR VPWR net3523 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11981_ clknet_leaf_14_clk _00789_ VGND VGND VPWR VPWR data_array.data0\[4\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_44_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1883 data_array.data0\[15\]\[15\] VGND VGND VPWR VPWR net3534 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13720_ clknet_leaf_214_clk _02349_ VGND VGND VPWR VPWR data_array.data1\[1\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_44_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1894 tag_array.tag1\[12\]\[10\] VGND VGND VPWR VPWR net3545 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_16_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10932_ net1014 net4144 net532 VGND VGND VPWR VPWR _02677_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_158_3406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_73 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13651_ clknet_leaf_35_clk _02280_ VGND VGND VPWR VPWR data_array.data1\[15\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_10863_ net1034 net2995 net520 VGND VGND VPWR VPWR _02608_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_175_3720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_175_3731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12602_ clknet_leaf_160_clk _01296_ VGND VGND VPWR VPWR tag_array.tag0\[0\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_71_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13582_ clknet_leaf_94_clk _02211_ VGND VGND VPWR VPWR data_array.data0\[9\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_10794_ net1848 net1054 net507 VGND VGND VPWR VPWR _02539_ sky130_fd_sc_hd__mux2_1
XFILLER_13_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12533_ clknet_leaf_99_clk _01227_ VGND VGND VPWR VPWR tag_array.tag1\[11\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_171_3639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12464_ clknet_leaf_213_clk _01158_ VGND VGND VPWR VPWR data_array.data1\[9\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14203_ clknet_leaf_2_clk _02832_ VGND VGND VPWR VPWR data_array.data0\[2\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
X_11415_ clknet_leaf_72_clk _00225_ VGND VGND VPWR VPWR data_array.data0\[0\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_12395_ clknet_leaf_206_clk _01089_ VGND VGND VPWR VPWR data_array.data0\[14\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_181_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14134_ clknet_leaf_6_clk _02763_ VGND VGND VPWR VPWR data_array.data0\[1\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_126_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11346_ net908 net3429 net797 VGND VGND VPWR VPWR _03089_ sky130_fd_sc_hd__mux2_1
XFILLER_152_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14065_ clknet_leaf_257_clk _02694_ VGND VGND VPWR VPWR data_array.data1\[6\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
X_11277_ net922 net3338 net682 VGND VGND VPWR VPWR _03020_ sky130_fd_sc_hd__mux2_1
XFILLER_165_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13016_ clknet_leaf_38_clk _01710_ VGND VGND VPWR VPWR data_array.data0\[3\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_10228_ net894 net3281 net356 VGND VGND VPWR VPWR _01975_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10159_ net910 net4379 net369 VGND VGND VPWR VPWR _01907_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13918_ clknet_leaf_24_clk _02547_ VGND VGND VPWR VPWR data_array.data1\[4\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_18_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13849_ clknet_leaf_253_clk _02478_ VGND VGND VPWR VPWR data_array.data1\[3\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_07370_ data_array.data0\[5\]\[57\] net1539 net1443 data_array.data0\[6\]\[57\] VGND
+ VGND VPWR VPWR _04618_ sky130_fd_sc_hd__a22o_1
XFILLER_176_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06321_ tag_array.tag0\[5\]\[12\] net1597 net1501 tag_array.tag0\[6\]\[12\] VGND
+ VGND VPWR VPWR _03664_ sky130_fd_sc_hd__a22o_1
XFILLER_31_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09040_ net2382 net866 net420 VGND VGND VPWR VPWR _00795_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_96_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06252_ _03600_ _03601_ VGND VGND VPWR VPWR _00151_ sky130_fd_sc_hd__or2_1
X_06183_ tag_array.valid1\[4\] net1366 net1273 tag_array.valid1\[7\] _03538_ VGND
+ VGND VPWR VPWR _03539_ sky130_fd_sc_hd__a221o_1
XFILLER_117_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold402 data_array.data0\[0\]\[36\] VGND VGND VPWR VPWR net2053 sky130_fd_sc_hd__dlygate4sd3_1
Xhold413 data_array.data0\[0\]\[27\] VGND VGND VPWR VPWR net2064 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold424 data_array.data1\[8\]\[60\] VGND VGND VPWR VPWR net2075 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold435 tag_array.tag1\[8\]\[24\] VGND VGND VPWR VPWR net2086 sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 data_array.data0\[8\]\[10\] VGND VGND VPWR VPWR net2097 sky130_fd_sc_hd__dlygate4sd3_1
Xhold457 data_array.data1\[8\]\[48\] VGND VGND VPWR VPWR net2108 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold468 data_array.data0\[2\]\[6\] VGND VGND VPWR VPWR net2119 sky130_fd_sc_hd__dlygate4sd3_1
X_09942_ net1060 net4343 net377 VGND VGND VPWR VPWR _01691_ sky130_fd_sc_hd__mux2_1
Xhold479 data_array.data1\[8\]\[1\] VGND VGND VPWR VPWR net2130 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout904 _05522_ VGND VGND VPWR VPWR net904 sky130_fd_sc_hd__clkbuf_2
XFILLER_98_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout915 _05518_ VGND VGND VPWR VPWR net915 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout926 _05512_ VGND VGND VPWR VPWR net926 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_70_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout937 net938 VGND VGND VPWR VPWR net937 sky130_fd_sc_hd__clkbuf_2
X_09873_ net976 net4328 net383 VGND VGND VPWR VPWR _01623_ sky130_fd_sc_hd__mux2_1
Xfanout948 _05500_ VGND VGND VPWR VPWR net948 sky130_fd_sc_hd__clkbuf_2
XFILLER_112_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout959 _05496_ VGND VGND VPWR VPWR net959 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1102 data_array.data1\[6\]\[40\] VGND VGND VPWR VPWR net2753 sky130_fd_sc_hd__dlygate4sd3_1
X_08824_ net1837 net949 net448 VGND VGND VPWR VPWR _00582_ sky130_fd_sc_hd__mux2_1
Xhold1113 tag_array.tag1\[1\]\[7\] VGND VGND VPWR VPWR net2764 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1124 tag_array.tag0\[11\]\[20\] VGND VGND VPWR VPWR net2775 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1135 data_array.data0\[4\]\[20\] VGND VGND VPWR VPWR net2786 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1146 data_array.data1\[1\]\[3\] VGND VGND VPWR VPWR net2797 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08755_ net702 net3228 net458 VGND VGND VPWR VPWR _00514_ sky130_fd_sc_hd__mux2_1
Xhold1157 tag_array.tag1\[5\]\[0\] VGND VGND VPWR VPWR net2808 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1168 data_array.data0\[15\]\[2\] VGND VGND VPWR VPWR net2819 sky130_fd_sc_hd__dlygate4sd3_1
X_05967_ data_array.rdata1\[45\] net829 net838 VGND VGND VPWR VPWR _03439_ sky130_fd_sc_hd__a21o_1
XFILLER_38_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1179 tag_array.tag0\[0\]\[18\] VGND VGND VPWR VPWR net2830 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07706_ data_array.data1\[12\]\[24\] net1395 net1301 data_array.data1\[15\]\[24\]
+ _04922_ VGND VGND VPWR VPWR _04923_ sky130_fd_sc_hd__a221o_1
X_08686_ net2042 net780 net482 VGND VGND VPWR VPWR _00445_ sky130_fd_sc_hd__mux2_1
X_05898_ data_array.rdata1\[22\] net829 net838 VGND VGND VPWR VPWR _03393_ sky130_fd_sc_hd__a21o_1
XFILLER_54_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07637_ net1214 _04855_ _04859_ net1166 VGND VGND VPWR VPWR _04861_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_68_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_105_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07568_ data_array.data1\[5\]\[11\] net1574 net1478 data_array.data1\[6\]\[11\] VGND
+ VGND VPWR VPWR _04798_ sky130_fd_sc_hd__a22o_1
XFILLER_179_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09307_ net750 net3545 net552 VGND VGND VPWR VPWR _01061_ sky130_fd_sc_hd__mux2_1
X_06519_ tag_array.tag1\[1\]\[5\] net1610 net1514 tag_array.tag1\[2\]\[5\] VGND VGND
+ VPWR VPWR _03844_ sky130_fd_sc_hd__a22o_1
XFILLER_16_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07499_ data_array.data1\[0\]\[5\] net1360 net1266 data_array.data1\[3\]\[5\] _04734_
+ VGND VGND VPWR VPWR _04735_ sky130_fd_sc_hd__a221o_1
XFILLER_70_59 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09238_ net727 net3189 net646 VGND VGND VPWR VPWR _00992_ sky130_fd_sc_hd__mux2_1
XFILLER_148_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09169_ net865 net3101 net570 VGND VGND VPWR VPWR _00923_ sky130_fd_sc_hd__mux2_1
XFILLER_163_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11200_ net975 net4017 net648 VGND VGND VPWR VPWR _02943_ sky130_fd_sc_hd__mux2_1
XFILLER_108_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12180_ clknet_leaf_163_clk _00988_ VGND VGND VPWR VPWR tag_array.tag0\[14\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11131_ net995 net4393 net548 VGND VGND VPWR VPWR _02874_ sky130_fd_sc_hd__mux2_1
XFILLER_135_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold980 data_array.data0\[12\]\[35\] VGND VGND VPWR VPWR net2631 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold991 tag_array.tag1\[12\]\[4\] VGND VGND VPWR VPWR net2642 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_168_3590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11062_ net2198 net1013 net333 VGND VGND VPWR VPWR _02805_ sky130_fd_sc_hd__mux2_1
XFILLER_49_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10013_ net1034 net2927 net562 VGND VGND VPWR VPWR _01762_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2370 data_array.data0\[5\]\[17\] VGND VGND VPWR VPWR net4021 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2381 data_array.data0\[12\]\[14\] VGND VGND VPWR VPWR net4032 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2392 data_array.data1\[5\]\[6\] VGND VGND VPWR VPWR net4043 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1680 data_array.data0\[11\]\[16\] VGND VGND VPWR VPWR net3331 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1691 data_array.data0\[6\]\[18\] VGND VGND VPWR VPWR net3342 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11964_ clknet_leaf_88_clk _00772_ VGND VGND VPWR VPWR data_array.data0\[4\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
X_13703_ clknet_leaf_193_clk _02332_ VGND VGND VPWR VPWR data_array.data1\[15\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
X_10915_ net1082 net4042 net532 VGND VGND VPWR VPWR _02660_ sky130_fd_sc_hd__mux2_1
X_11895_ clknet_leaf_90_clk _00703_ VGND VGND VPWR VPWR data_array.data0\[5\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_17_Left_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13634_ clknet_leaf_54_clk _02263_ VGND VGND VPWR VPWR data_array.data0\[9\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
X_10846_ net1100 net2634 net515 VGND VGND VPWR VPWR _02591_ sky130_fd_sc_hd__mux2_1
XFILLER_158_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13565_ clknet_leaf_123_clk _02194_ VGND VGND VPWR VPWR data_array.data1\[0\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10777_ net865 net3859 net494 VGND VGND VPWR VPWR _02522_ sky130_fd_sc_hd__mux2_1
XFILLER_8_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12516_ clknet_leaf_176_clk _01210_ VGND VGND VPWR VPWR lru_array.lru_mem\[1\] sky130_fd_sc_hd__dfxtp_1
X_13496_ clknet_leaf_35_clk _02125_ VGND VGND VPWR VPWR tag_array.dirty1\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_173_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12447_ clknet_leaf_178_clk _01141_ VGND VGND VPWR VPWR lru_array.lru_mem\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_154_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12378_ clknet_leaf_119_clk _00056_ VGND VGND VPWR VPWR data_array.rdata0\[60\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_26_Left_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14117_ clknet_leaf_52_clk _02746_ VGND VGND VPWR VPWR data_array.data0\[1\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_11329_ net978 net3738 net802 VGND VGND VPWR VPWR _03072_ sky130_fd_sc_hd__mux2_1
XFILLER_4_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14048_ clknet_leaf_91_clk _02677_ VGND VGND VPWR VPWR data_array.data1\[6\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_79_250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_892 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06870_ data_array.data0\[8\]\[12\] net1406 net1312 data_array.data0\[11\]\[12\]
+ _04162_ VGND VGND VPWR VPWR _04163_ sky130_fd_sc_hd__a221o_1
XFILLER_67_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05821_ _03334_ _03335_ _03336_ _03337_ VGND VGND VPWR VPWR _03338_ sky130_fd_sc_hd__or4_1
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_89_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08540_ net1715 net540 VGND VGND VPWR VPWR _00308_ sky130_fd_sc_hd__nand2b_1
X_05752_ net25 fsm.tag_out1\[24\] VGND VGND VPWR VPWR _03269_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_35_Left_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08471_ net1626 net1279 VGND VGND VPWR VPWR _05550_ sky130_fd_sc_hd__nand2_1
X_05683_ net22 fsm.tag_out0\[22\] VGND VGND VPWR VPWR _03200_ sky130_fd_sc_hd__and2b_1
X_07422_ data_array.data0\[4\]\[62\] net1412 net1318 data_array.data0\[7\]\[62\] _04664_
+ VGND VGND VPWR VPWR _04665_ sky130_fd_sc_hd__a221o_1
XFILLER_23_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07353_ data_array.data0\[13\]\[56\] net1531 net1435 data_array.data0\[14\]\[56\]
+ VGND VGND VPWR VPWR _04602_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_63_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06304_ tag_array.tag0\[0\]\[10\] net1404 net1310 tag_array.tag0\[3\]\[10\] _03648_
+ VGND VGND VPWR VPWR _03649_ sky130_fd_sc_hd__a221o_1
XFILLER_31_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07284_ net1204 _04533_ _04537_ net1630 VGND VGND VPWR VPWR _04540_ sky130_fd_sc_hd__a22o_1
XFILLER_176_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09023_ net1984 net932 net424 VGND VGND VPWR VPWR _00778_ sky130_fd_sc_hd__mux2_1
X_06235_ tag_array.tag0\[13\]\[4\] net1564 net1468 tag_array.tag0\[14\]\[4\] VGND
+ VGND VPWR VPWR _03586_ sky130_fd_sc_hd__a22o_1
XFILLER_156_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1051 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold210 data_array.data1\[1\]\[35\] VGND VGND VPWR VPWR net1861 sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 data_array.data1\[1\]\[10\] VGND VGND VPWR VPWR net1872 sky130_fd_sc_hd__dlygate4sd3_1
X_06166_ net28 net29 VGND VGND VPWR VPWR _03523_ sky130_fd_sc_hd__nand2_1
Xhold232 data_array.data0\[8\]\[22\] VGND VGND VPWR VPWR net1883 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold243 data_array.data0\[11\]\[15\] VGND VGND VPWR VPWR net1894 sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 data_array.data0\[0\]\[23\] VGND VGND VPWR VPWR net1905 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06097_ data_array.rdata0\[12\] net1141 net1119 data_array.rdata1\[12\] VGND VGND
+ VPWR VPWR net266 sky130_fd_sc_hd__a22o_1
Xhold265 data_array.data0\[4\]\[8\] VGND VGND VPWR VPWR net1916 sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 data_array.data0\[1\]\[6\] VGND VGND VPWR VPWR net1927 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold287 data_array.data0\[1\]\[22\] VGND VGND VPWR VPWR net1938 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout701 _05411_ VGND VGND VPWR VPWR net701 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold298 data_array.data0\[0\]\[51\] VGND VGND VPWR VPWR net1949 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout712 net713 VGND VGND VPWR VPWR net712 sky130_fd_sc_hd__clkbuf_2
X_09925_ net708 net2622 net604 VGND VGND VPWR VPWR _01675_ sky130_fd_sc_hd__mux2_1
Xfanout723 _05399_ VGND VGND VPWR VPWR net723 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout734 net735 VGND VGND VPWR VPWR net734 sky130_fd_sc_hd__clkbuf_2
Xfanout745 _05389_ VGND VGND VPWR VPWR net745 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout756 _05383_ VGND VGND VPWR VPWR net756 sky130_fd_sc_hd__clkbuf_2
X_09856_ net1046 net3626 net380 VGND VGND VPWR VPWR _01606_ sky130_fd_sc_hd__mux2_1
Xfanout767 _05377_ VGND VGND VPWR VPWR net767 sky130_fd_sc_hd__buf_1
Xfanout778 net779 VGND VGND VPWR VPWR net778 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_146_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout789 net790 VGND VGND VPWR VPWR net789 sky130_fd_sc_hd__clkbuf_2
X_08807_ net4310 net1019 net444 VGND VGND VPWR VPWR _00565_ sky130_fd_sc_hd__mux2_1
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09787_ net1061 net2469 net392 VGND VGND VPWR VPWR _01538_ sky130_fd_sc_hd__mux2_1
X_06999_ net1221 _04275_ _04279_ net1172 VGND VGND VPWR VPWR _04281_ sky130_fd_sc_hd__a22o_1
XFILLER_61_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08738_ net772 net4173 net463 VGND VGND VPWR VPWR _00497_ sky130_fd_sc_hd__mux2_1
XFILLER_22_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08669_ net746 net3183 net499 VGND VGND VPWR VPWR _00428_ sky130_fd_sc_hd__mux2_1
X_10700_ net2891 net918 net484 VGND VGND VPWR VPWR _02445_ sky130_fd_sc_hd__mux2_1
XFILLER_41_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11680_ clknet_leaf_100_clk _00488_ VGND VGND VPWR VPWR tag_array.tag1\[1\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_120_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10631_ net2110 net937 net471 VGND VGND VPWR VPWR _02376_ sky130_fd_sc_hd__mux2_1
XFILLER_14_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13350_ clknet_leaf_54_clk _01980_ VGND VGND VPWR VPWR data_array.data0\[10\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
X_10562_ net958 net3317 net461 VGND VGND VPWR VPWR _02307_ sky130_fd_sc_hd__mux2_1
XFILLER_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12301_ clknet_leaf_137_clk _01059_ VGND VGND VPWR VPWR tag_array.tag1\[12\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_13281_ clknet_leaf_223_clk _01911_ VGND VGND VPWR VPWR data_array.data0\[11\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_20_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10493_ net972 net3749 net344 VGND VGND VPWR VPWR _02238_ sky130_fd_sc_hd__mux2_1
XFILLER_182_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12232_ clknet_leaf_182_clk _00161_ VGND VGND VPWR VPWR fsm.tag_out1\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_931 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12163_ clknet_leaf_171_clk _00971_ VGND VGND VPWR VPWR tag_array.tag0\[13\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_123_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_166_3549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11114_ net1063 net3922 net550 VGND VGND VPWR VPWR _02857_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12094_ clknet_leaf_122_clk _00902_ VGND VGND VPWR VPWR data_array.data1\[14\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_183_3874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11045_ net3028 net1081 net335 VGND VGND VPWR VPWR _02788_ sky130_fd_sc_hd__mux2_1
XFILLER_118_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12996_ clknet_leaf_45_clk _01690_ VGND VGND VPWR VPWR data_array.data0\[3\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11947_ clknet_leaf_228_clk _00755_ VGND VGND VPWR VPWR data_array.data0\[4\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11878_ clknet_leaf_223_clk _00686_ VGND VGND VPWR VPWR data_array.data0\[5\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_13617_ clknet_leaf_93_clk _02246_ VGND VGND VPWR VPWR data_array.data0\[9\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10829_ net2231 net915 net508 VGND VGND VPWR VPWR _02574_ sky130_fd_sc_hd__mux2_1
XFILLER_32_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13548_ clknet_leaf_26_clk _02177_ VGND VGND VPWR VPWR data_array.data1\[0\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_173_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13479_ clknet_leaf_108_clk _02109_ VGND VGND VPWR VPWR tag_array.tag0\[15\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06020_ data_array.rdata0\[63\] net849 net1144 VGND VGND VPWR VPWR _03474_ sky130_fd_sc_hd__o21a_1
Xoutput304 net304 VGND VGND VPWR VPWR mem_wdata[47] sky130_fd_sc_hd__buf_2
XFILLER_161_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput315 net315 VGND VGND VPWR VPWR mem_wdata[57] sky130_fd_sc_hd__buf_2
Xoutput326 net326 VGND VGND VPWR VPWR mem_wdata[9] sky130_fd_sc_hd__buf_2
XFILLER_113_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07971_ data_array.data1\[5\]\[48\] net1583 net1487 data_array.data1\[6\]\[48\] VGND
+ VGND VPWR VPWR _05164_ sky130_fd_sc_hd__a22o_1
XFILLER_99_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09710_ net748 net3750 net609 VGND VGND VPWR VPWR _01462_ sky130_fd_sc_hd__mux2_1
X_06922_ net1174 _04205_ _04209_ net1220 VGND VGND VPWR VPWR _04211_ sky130_fd_sc_hd__a22o_1
X_09641_ net723 net2831 net616 VGND VGND VPWR VPWR _01393_ sky130_fd_sc_hd__mux2_1
X_06853_ data_array.data0\[1\]\[10\] net1601 net1505 data_array.data0\[2\]\[10\] VGND
+ VGND VPWR VPWR _04148_ sky130_fd_sc_hd__a22o_1
X_05804_ _03195_ _03201_ VGND VGND VPWR VPWR _03321_ sky130_fd_sc_hd__or2_1
XFILLER_83_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09572_ net1061 net3108 net400 VGND VGND VPWR VPWR _01324_ sky130_fd_sc_hd__mux2_1
X_06784_ data_array.data0\[4\]\[4\] net1391 net1297 data_array.data0\[7\]\[4\] _04084_
+ VGND VGND VPWR VPWR _04085_ sky130_fd_sc_hd__a221o_1
XFILLER_83_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_141_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08523_ net1712 net597 VGND VGND VPWR VPWR _00302_ sky130_fd_sc_hd__nand2b_1
XFILLER_42_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05735_ net15 fsm.tag_out1\[15\] VGND VGND VPWR VPWR _03252_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_65_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08454_ net155 net90 net1648 VGND VGND VPWR VPWR _05539_ sky130_fd_sc_hd__mux2_1
X_05666_ net6 fsm.tag_out0\[7\] VGND VGND VPWR VPWR _03183_ sky130_fd_sc_hd__and2b_1
XFILLER_23_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07405_ net1635 _04643_ _04647_ net1209 VGND VGND VPWR VPWR _04650_ sky130_fd_sc_hd__a22o_1
X_08385_ net129 net64 net1643 VGND VGND VPWR VPWR _05493_ sky130_fd_sc_hd__mux2_1
X_07336_ data_array.data0\[12\]\[54\] net1356 net1262 data_array.data0\[15\]\[54\]
+ _04586_ VGND VGND VPWR VPWR _04587_ sky130_fd_sc_hd__a221o_1
XFILLER_137_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07267_ data_array.data0\[5\]\[48\] net1578 net1482 data_array.data0\[6\]\[48\] VGND
+ VGND VPWR VPWR _04524_ sky130_fd_sc_hd__a22o_1
XFILLER_164_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09006_ net2274 net1003 net420 VGND VGND VPWR VPWR _00761_ sky130_fd_sc_hd__mux2_1
X_06218_ net1181 _03565_ _03569_ net1229 VGND VGND VPWR VPWR _03571_ sky130_fd_sc_hd__a22o_1
XFILLER_164_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07198_ _04460_ _04461_ VGND VGND VPWR VPWR _00035_ sky130_fd_sc_hd__or2_1
XFILLER_145_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06149_ net28 net29 VGND VGND VPWR VPWR _03506_ sky130_fd_sc_hd__and2b_4
XFILLER_104_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_6_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1507 net1516 VGND VGND VPWR VPWR net1507 sky130_fd_sc_hd__clkbuf_4
Xfanout1518 _03510_ VGND VGND VPWR VPWR net1518 sky130_fd_sc_hd__buf_4
Xfanout520 net522 VGND VGND VPWR VPWR net520 sky130_fd_sc_hd__clkbuf_8
Xfanout1529 net1530 VGND VGND VPWR VPWR net1529 sky130_fd_sc_hd__clkbuf_2
Xfanout531 net534 VGND VGND VPWR VPWR net531 sky130_fd_sc_hd__clkbuf_8
Xfanout542 net547 VGND VGND VPWR VPWR net542 sky130_fd_sc_hd__clkbuf_4
X_09908_ net777 net4333 net602 VGND VGND VPWR VPWR _01658_ sky130_fd_sc_hd__mux2_1
Xfanout553 _05594_ VGND VGND VPWR VPWR net553 sky130_fd_sc_hd__clkbuf_4
Xfanout564 net565 VGND VGND VPWR VPWR net564 sky130_fd_sc_hd__buf_4
Xfanout575 _05592_ VGND VGND VPWR VPWR net575 sky130_fd_sc_hd__buf_4
Xfanout586 net590 VGND VGND VPWR VPWR net586 sky130_fd_sc_hd__clkbuf_8
X_09839_ _05414_ _05558_ VGND VGND VPWR VPWR _03126_ sky130_fd_sc_hd__or2_1
Xfanout597 net598 VGND VGND VPWR VPWR net597 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_161_3457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12850_ clknet_leaf_16_clk _01544_ VGND VGND VPWR VPWR data_array.data0\[12\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_122_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_122_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ clknet_leaf_48_clk _00609_ VGND VGND VPWR VPWR data_array.data0\[7\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12781_ clknet_leaf_177_clk _01475_ VGND VGND VPWR VPWR tag_array.tag0\[6\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11732_ clknet_leaf_143_clk _00540_ VGND VGND VPWR VPWR tag_array.tag0\[9\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_25_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ clknet_leaf_256_clk _03074_ VGND VGND VPWR VPWR data_array.data1\[7\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
X_11663_ clknet_leaf_194_clk _00471_ VGND VGND VPWR VPWR tag_array.tag1\[1\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_153_Right_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13402_ clknet_leaf_25_clk _02032_ VGND VGND VPWR VPWR data_array.data1\[8\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_10614_ net1762 net1005 net468 VGND VGND VPWR VPWR _02359_ sky130_fd_sc_hd__mux2_1
X_14382_ clknet_leaf_265_clk _03005_ VGND VGND VPWR VPWR data_array.data1\[10\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_155_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11594_ clknet_leaf_102_clk _00402_ VGND VGND VPWR VPWR tag_array.tag1\[4\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_13333_ clknet_leaf_93_clk _01963_ VGND VGND VPWR VPWR data_array.data0\[10\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
X_10545_ net1024 net2991 net454 VGND VGND VPWR VPWR _02290_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_130_clk clknet_5_30__leaf_clk VGND VGND VPWR VPWR clknet_leaf_130_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13264_ clknet_leaf_223_clk _01894_ VGND VGND VPWR VPWR data_array.data0\[11\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_155_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10476_ net1043 net2931 net344 VGND VGND VPWR VPWR _02221_ sky130_fd_sc_hd__mux2_1
X_12215_ clknet_leaf_184_clk _00145_ VGND VGND VPWR VPWR fsm.tag_out0\[22\] sky130_fd_sc_hd__dfxtp_2
X_13195_ clknet_leaf_257_clk _00089_ VGND VGND VPWR VPWR data_array.rdata1\[32\] sky130_fd_sc_hd__dfxtp_1
X_12146_ clknet_leaf_171_clk _00954_ VGND VGND VPWR VPWR tag_array.tag0\[13\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_111_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12077_ clknet_leaf_204_clk _00885_ VGND VGND VPWR VPWR data_array.data1\[14\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_49_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11028_ net1999 net888 net337 VGND VGND VPWR VPWR _02772_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_197_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_197_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12979_ clknet_leaf_106_clk _01673_ VGND VGND VPWR VPWR tag_array.tag0\[4\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_43_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_16 _03154_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_120_Right_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_27 _05411_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_38 net470 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08170_ lru_array.lru_mem\[4\] net1371 net1277 lru_array.lru_mem\[7\] _05344_ VGND
+ VGND VPWR VPWR _05345_ sky130_fd_sc_hd__a221o_1
XANTENNA_49 net666 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07121_ _04390_ _04391_ VGND VGND VPWR VPWR _00027_ sky130_fd_sc_hd__or2_1
XFILLER_118_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_121_clk clknet_5_27__leaf_clk VGND VGND VPWR VPWR clknet_leaf_121_clk
+ sky130_fd_sc_hd__clkbuf_8
X_07052_ data_array.data0\[0\]\[28\] net1350 net1256 data_array.data0\[3\]\[28\] _04328_
+ VGND VGND VPWR VPWR _04329_ sky130_fd_sc_hd__a221o_1
XFILLER_146_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06003_ data_array.rdata1\[57\] net830 net839 VGND VGND VPWR VPWR _03463_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_58_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput167 net167 VGND VGND VPWR VPWR cpu_rdata[11] sky130_fd_sc_hd__buf_6
Xoutput178 net178 VGND VGND VPWR VPWR cpu_rdata[21] sky130_fd_sc_hd__clkbuf_4
Xoutput189 net189 VGND VGND VPWR VPWR cpu_rdata[31] sky130_fd_sc_hd__buf_6
XFILLER_87_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2903 tag_array.tag0\[13\]\[19\] VGND VGND VPWR VPWR net4554 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2914 data_array.data1\[6\]\[61\] VGND VGND VPWR VPWR net4565 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2925 data_array.data1\[5\]\[32\] VGND VGND VPWR VPWR net4576 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2936 data_array.data0\[5\]\[20\] VGND VGND VPWR VPWR net4587 sky130_fd_sc_hd__dlygate4sd3_1
X_07954_ data_array.data1\[0\]\[46\] net1333 net1239 data_array.data1\[3\]\[46\] _05148_
+ VGND VGND VPWR VPWR _05149_ sky130_fd_sc_hd__a221o_1
Xhold2947 tag_array.tag0\[7\]\[16\] VGND VGND VPWR VPWR net4598 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_143_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2958 data_array.data1\[5\]\[12\] VGND VGND VPWR VPWR net4609 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_143_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06905_ data_array.data0\[4\]\[15\] net1390 net1296 data_array.data0\[7\]\[15\] _04194_
+ VGND VGND VPWR VPWR _04195_ sky130_fd_sc_hd__a221o_1
Xhold2969 data_array.data1\[6\]\[12\] VGND VGND VPWR VPWR net4620 sky130_fd_sc_hd__dlygate4sd3_1
X_07885_ data_array.data1\[9\]\[40\] net1605 net1509 data_array.data1\[10\]\[40\]
+ VGND VGND VPWR VPWR _05086_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_188_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_188_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_29_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09624_ net794 net3011 net616 VGND VGND VPWR VPWR _01376_ sky130_fd_sc_hd__mux2_1
XFILLER_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06836_ data_array.data0\[9\]\[9\] net1580 net1484 data_array.data0\[10\]\[9\] VGND
+ VGND VPWR VPWR _04132_ sky130_fd_sc_hd__a22o_1
XFILLER_83_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09555_ net708 net2511 net620 VGND VGND VPWR VPWR _01308_ sky130_fd_sc_hd__mux2_1
X_06767_ net1190 _04063_ _04067_ net1616 VGND VGND VPWR VPWR _04070_ sky130_fd_sc_hd__a22o_1
XFILLER_43_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08506_ _03511_ _03527_ VGND VGND VPWR VPWR _05574_ sky130_fd_sc_hd__nor2_1
XFILLER_102_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05718_ _03232_ _03233_ _03234_ VGND VGND VPWR VPWR _03235_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_80_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09486_ net784 net2293 net624 VGND VGND VPWR VPWR _01239_ sky130_fd_sc_hd__mux2_1
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06698_ tag_array.tag1\[12\]\[21\] net1404 net1310 tag_array.tag1\[15\]\[21\] _04006_
+ VGND VGND VPWR VPWR _04007_ sky130_fd_sc_hd__a221o_1
XFILLER_178_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08437_ net1125 _05527_ VGND VGND VPWR VPWR _05528_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_22_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05649_ _03164_ _03165_ _03163_ VGND VGND VPWR VPWR _03166_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_22_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08368_ net1128 _05481_ VGND VGND VPWR VPWR _05482_ sky130_fd_sc_hd__and2_1
XFILLER_137_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07319_ _04570_ _04571_ VGND VGND VPWR VPWR _00047_ sky130_fd_sc_hd__or2_1
XFILLER_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08299_ net1124 _05435_ VGND VGND VPWR VPWR _05436_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_112_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_112_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_137_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10330_ net780 net3828 net591 VGND VGND VPWR VPWR _02077_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_115_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10261_ net699 net2905 net596 VGND VGND VPWR VPWR _02008_ sky130_fd_sc_hd__mux2_1
XFILLER_79_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12000_ clknet_leaf_112_clk _00808_ VGND VGND VPWR VPWR data_array.data0\[6\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10192_ net1037 net4068 net358 VGND VGND VPWR VPWR _01939_ sky130_fd_sc_hd__mux2_1
XFILLER_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1304 net1305 VGND VGND VPWR VPWR net1304 sky130_fd_sc_hd__clkbuf_4
Xfanout1315 net1328 VGND VGND VPWR VPWR net1315 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_180_3811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1326 net1327 VGND VGND VPWR VPWR net1326 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_180_3822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1337 net1338 VGND VGND VPWR VPWR net1337 sky130_fd_sc_hd__clkbuf_4
Xfanout1348 net1352 VGND VGND VPWR VPWR net1348 sky130_fd_sc_hd__buf_2
Xfanout350 net351 VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__clkbuf_8
Xfanout361 _03129_ VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__buf_4
Xfanout1359 net1360 VGND VGND VPWR VPWR net1359 sky130_fd_sc_hd__clkbuf_4
XFILLER_93_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout372 net373 VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__buf_4
XFILLER_143_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout383 net384 VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__buf_4
X_13951_ clknet_leaf_21_clk _02580_ VGND VGND VPWR VPWR data_array.data1\[4\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_179_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_179_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_115_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout394 net395 VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__clkbuf_8
XFILLER_86_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12902_ clknet_leaf_0_clk _01596_ VGND VGND VPWR VPWR data_array.data0\[13\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13882_ clknet_leaf_246_clk _02511_ VGND VGND VPWR VPWR data_array.data1\[3\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12833_ clknet_leaf_261_clk _01527_ VGND VGND VPWR VPWR data_array.data0\[12\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_178_3773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ clknet_leaf_143_clk _01458_ VGND VGND VPWR VPWR tag_array.tag0\[6\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_178_3784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11715_ clknet_leaf_179_clk _00523_ VGND VGND VPWR VPWR tag_array.tag0\[9\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_12695_ clknet_leaf_147_clk _01389_ VGND VGND VPWR VPWR tag_array.tag0\[8\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_159_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14434_ clknet_leaf_18_clk _03057_ VGND VGND VPWR VPWR data_array.data1\[7\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_11646_ clknet_leaf_99_clk _00454_ VGND VGND VPWR VPWR tag_array.tag1\[2\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput14 cpu_addr[21] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_2
XFILLER_174_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14365_ clknet_leaf_70_clk _02988_ VGND VGND VPWR VPWR data_array.data1\[10\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput25 cpu_addr[31] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__buf_1
X_11577_ clknet_leaf_189_clk _00385_ VGND VGND VPWR VPWR tag_array.tag1\[5\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput36 cpu_wdata[11] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_103_clk clknet_5_24__leaf_clk VGND VGND VPWR VPWR clknet_leaf_103_clk
+ sky130_fd_sc_hd__clkbuf_8
Xinput47 cpu_wdata[21] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_1
X_13316_ clknet_leaf_0_clk _01946_ VGND VGND VPWR VPWR data_array.data0\[10\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput58 cpu_wdata[31] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_1
X_10528_ net1094 net4185 net461 VGND VGND VPWR VPWR _02273_ sky130_fd_sc_hd__mux2_1
Xinput69 cpu_wdata[41] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__clkbuf_1
Xhold809 data_array.data1\[14\]\[10\] VGND VGND VPWR VPWR net2460 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_824 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14296_ clknet_leaf_213_clk _02925_ VGND VGND VPWR VPWR data_array.data1\[11\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_109_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13247_ clknet_leaf_126_clk _01877_ VGND VGND VPWR VPWR data_array.data0\[11\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_10459_ net1109 net2869 net346 VGND VGND VPWR VPWR _02204_ sky130_fd_sc_hd__mux2_1
XFILLER_184_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13178_ clknet_leaf_65_clk _00070_ VGND VGND VPWR VPWR data_array.rdata1\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_69_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12129_ clknet_leaf_163_clk _00937_ VGND VGND VPWR VPWR tag_array.tag0\[12\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_36_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1509 tag_array.tag0\[5\]\[0\] VGND VGND VPWR VPWR net3160 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_42_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07670_ net1185 _04885_ _04889_ net1233 VGND VGND VPWR VPWR _04891_ sky130_fd_sc_hd__a22o_1
XFILLER_37_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06621_ tag_array.tag1\[12\]\[14\] net1368 net1274 tag_array.tag1\[15\]\[14\] _03936_
+ VGND VGND VPWR VPWR _03937_ sky130_fd_sc_hd__a221o_1
XFILLER_53_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09340_ net1043 net3966 net404 VGND VGND VPWR VPWR _01093_ sky130_fd_sc_hd__mux2_1
X_06552_ tag_array.tag1\[5\]\[8\] net1609 net1513 tag_array.tag1\[6\]\[8\] VGND VGND
+ VPWR VPWR _03874_ sky130_fd_sc_hd__a22o_1
XFILLER_178_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09271_ net695 net2123 net571 VGND VGND VPWR VPWR _01025_ sky130_fd_sc_hd__mux2_1
XFILLER_61_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06483_ _03810_ _03811_ VGND VGND VPWR VPWR _00167_ sky130_fd_sc_hd__or2_2
XFILLER_20_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08222_ fsm.tag_out1\[9\] net817 net809 fsm.tag_out0\[9\] _05382_ VGND VGND VPWR
+ VPWR _05383_ sky130_fd_sc_hd__a221o_2
XFILLER_159_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08153_ net1193 _05323_ _05327_ net1619 VGND VGND VPWR VPWR _05330_ sky130_fd_sc_hd__a22o_1
XFILLER_174_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07104_ data_array.data0\[9\]\[33\] net1585 net1489 data_array.data0\[10\]\[33\]
+ VGND VGND VPWR VPWR _04376_ sky130_fd_sc_hd__a22o_1
XFILLER_180_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload230 clknet_leaf_128_clk VGND VGND VPWR VPWR clkload230/Y sky130_fd_sc_hd__inv_8
X_08084_ data_array.data1\[12\]\[58\] net1359 net1265 data_array.data1\[15\]\[58\]
+ _05266_ VGND VGND VPWR VPWR _05267_ sky130_fd_sc_hd__a221o_1
Xclkload241 clknet_leaf_138_clk VGND VGND VPWR VPWR clkload241/Y sky130_fd_sc_hd__inv_8
X_07035_ data_array.data0\[8\]\[27\] net1367 net1273 data_array.data0\[11\]\[27\]
+ _04312_ VGND VGND VPWR VPWR _04313_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_77_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2700 data_array.data0\[7\]\[27\] VGND VGND VPWR VPWR net4351 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_73_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2711 data_array.data1\[11\]\[33\] VGND VGND VPWR VPWR net4362 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_110_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2722 tag_array.tag1\[9\]\[21\] VGND VGND VPWR VPWR net4373 sky130_fd_sc_hd__dlygate4sd3_1
X_08986_ net1988 net1080 net424 VGND VGND VPWR VPWR _00741_ sky130_fd_sc_hd__mux2_1
Xhold2733 data_array.data0\[11\]\[1\] VGND VGND VPWR VPWR net4384 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_110_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2744 data_array.data1\[14\]\[56\] VGND VGND VPWR VPWR net4395 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2755 data_array.data1\[10\]\[41\] VGND VGND VPWR VPWR net4406 sky130_fd_sc_hd__dlygate4sd3_1
X_07937_ data_array.data1\[12\]\[45\] net1350 net1256 data_array.data1\[15\]\[45\]
+ _05132_ VGND VGND VPWR VPWR _05133_ sky130_fd_sc_hd__a221o_1
Xhold2766 tag_array.tag0\[1\]\[9\] VGND VGND VPWR VPWR net4417 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2777 data_array.data0\[15\]\[50\] VGND VGND VPWR VPWR net4428 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2788 tag_array.tag1\[9\]\[1\] VGND VGND VPWR VPWR net4439 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2799 tag_array.tag1\[9\]\[19\] VGND VGND VPWR VPWR net4450 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07868_ net1228 _05065_ _05069_ net1180 VGND VGND VPWR VPWR _05071_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_27_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09607_ net920 net3698 net398 VGND VGND VPWR VPWR _01359_ sky130_fd_sc_hd__mux2_1
X_06819_ data_array.data0\[12\]\[7\] net1411 net1317 data_array.data0\[15\]\[7\] _04116_
+ VGND VGND VPWR VPWR _04117_ sky130_fd_sc_hd__a221o_1
X_07799_ data_array.data1\[5\]\[32\] net1520 net1424 data_array.data1\[6\]\[32\] VGND
+ VGND VPWR VPWR _05008_ sky130_fd_sc_hd__a22o_1
X_09538_ net776 net4202 net618 VGND VGND VPWR VPWR _01291_ sky130_fd_sc_hd__mux2_1
XFILLER_25_985 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09469_ net751 net2621 net659 VGND VGND VPWR VPWR _01222_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_156_3356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11500_ clknet_leaf_157_clk _00308_ VGND VGND VPWR VPWR tag_array.valid0\[15\] sky130_fd_sc_hd__dfxtp_1
X_12480_ clknet_leaf_265_clk _01174_ VGND VGND VPWR VPWR data_array.data1\[9\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11431_ clknet_leaf_126_clk _00241_ VGND VGND VPWR VPWR data_array.data0\[0\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_117_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14150_ clknet_leaf_109_clk _02779_ VGND VGND VPWR VPWR data_array.data0\[1\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11362_ net1648 net4468 net592 VGND VGND VPWR VPWR _03105_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_134_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13101_ clknet_leaf_208_clk _01795_ VGND VGND VPWR VPWR data_array.data1\[13\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
X_10313_ net1835 net910 net634 VGND VGND VPWR VPWR _02060_ sky130_fd_sc_hd__mux2_1
XFILLER_98_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14081_ clknet_leaf_249_clk _02710_ VGND VGND VPWR VPWR data_array.data1\[6\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11293_ net859 net3371 net678 VGND VGND VPWR VPWR _03036_ sky130_fd_sc_hd__mux2_1
X_13032_ clknet_leaf_91_clk _01726_ VGND VGND VPWR VPWR data_array.data0\[3\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_79_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10244_ net768 net3632 net595 VGND VGND VPWR VPWR _01991_ sky130_fd_sc_hd__mux2_1
Xfanout1101 _05424_ VGND VGND VPWR VPWR net1101 sky130_fd_sc_hd__buf_1
XFILLER_3_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1112 net1113 VGND VGND VPWR VPWR net1112 sky130_fd_sc_hd__buf_4
X_10175_ net1105 net4621 net354 VGND VGND VPWR VPWR _01922_ sky130_fd_sc_hd__mux2_1
XFILLER_79_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1123 net1124 VGND VGND VPWR VPWR net1123 sky130_fd_sc_hd__buf_4
Xfanout1134 net1135 VGND VGND VPWR VPWR net1134 sky130_fd_sc_hd__buf_4
XFILLER_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1145 net1146 VGND VGND VPWR VPWR net1145 sky130_fd_sc_hd__clkbuf_4
XFILLER_93_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1156 net1157 VGND VGND VPWR VPWR net1156 sky130_fd_sc_hd__buf_4
Xfanout1167 net1175 VGND VGND VPWR VPWR net1167 sky130_fd_sc_hd__clkbuf_4
Xfanout1178 net1180 VGND VGND VPWR VPWR net1178 sky130_fd_sc_hd__buf_4
XFILLER_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1189 net1191 VGND VGND VPWR VPWR net1189 sky130_fd_sc_hd__clkbuf_2
XFILLER_75_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13934_ clknet_leaf_74_clk _02563_ VGND VGND VPWR VPWR data_array.data1\[4\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13865_ clknet_leaf_73_clk _02494_ VGND VGND VPWR VPWR data_array.data1\[3\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_395 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12816_ clknet_leaf_127_clk _01510_ VGND VGND VPWR VPWR tag_array.tag1\[0\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_13796_ clknet_leaf_234_clk _02425_ VGND VGND VPWR VPWR data_array.data1\[2\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_43_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12747_ clknet_leaf_165_clk _01441_ VGND VGND VPWR VPWR tag_array.tag0\[5\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_176_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12678_ clknet_leaf_110_clk _01372_ VGND VGND VPWR VPWR data_array.data0\[15\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_13_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14417_ clknet_leaf_266_clk _03040_ VGND VGND VPWR VPWR data_array.data1\[7\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11629_ clknet_leaf_232_clk _00437_ VGND VGND VPWR VPWR tag_array.tag1\[3\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14348_ clknet_leaf_184_clk _00188_ _00193_ VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__dfrtp_1
XFILLER_128_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold606 data_array.data1\[0\]\[16\] VGND VGND VPWR VPWR net2257 sky130_fd_sc_hd__dlygate4sd3_1
Xhold617 data_array.data0\[8\]\[6\] VGND VGND VPWR VPWR net2268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold628 tag_array.tag1\[1\]\[16\] VGND VGND VPWR VPWR net2279 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14279_ clknet_leaf_193_clk _02908_ VGND VGND VPWR VPWR data_array.data1\[12\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold639 tag_array.tag1\[2\]\[24\] VGND VGND VPWR VPWR net2290 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_94_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2007 data_array.data0\[2\]\[30\] VGND VGND VPWR VPWR net3658 sky130_fd_sc_hd__dlygate4sd3_1
X_08840_ net2079 net885 net443 VGND VGND VPWR VPWR _00598_ sky130_fd_sc_hd__mux2_1
Xhold2018 data_array.data1\[11\]\[10\] VGND VGND VPWR VPWR net3669 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2029 tag_array.tag1\[1\]\[9\] VGND VGND VPWR VPWR net3680 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1306 data_array.data1\[5\]\[58\] VGND VGND VPWR VPWR net2957 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1317 tag_array.tag1\[6\]\[2\] VGND VGND VPWR VPWR net2968 sky130_fd_sc_hd__dlygate4sd3_1
X_08771_ net739 net4122 net452 VGND VGND VPWR VPWR _00530_ sky130_fd_sc_hd__mux2_1
Xhold1328 data_array.data1\[3\]\[40\] VGND VGND VPWR VPWR net2979 sky130_fd_sc_hd__dlygate4sd3_1
X_05983_ net144 net1150 _03448_ _03449_ VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__a22o_1
XFILLER_85_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1339 tag_array.tag1\[9\]\[5\] VGND VGND VPWR VPWR net2990 sky130_fd_sc_hd__dlygate4sd3_1
X_07722_ data_array.data1\[5\]\[25\] net1519 net1423 data_array.data1\[6\]\[25\] VGND
+ VGND VPWR VPWR _04938_ sky130_fd_sc_hd__a22o_1
XFILLER_66_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07653_ data_array.data1\[4\]\[19\] net1394 net1300 data_array.data1\[7\]\[19\] _04874_
+ VGND VGND VPWR VPWR _04875_ sky130_fd_sc_hd__a221o_1
XFILLER_81_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06604_ _03920_ _03921_ VGND VGND VPWR VPWR _00159_ sky130_fd_sc_hd__or2_1
X_07584_ data_array.data1\[13\]\[13\] net1551 net1455 data_array.data1\[14\]\[13\]
+ VGND VGND VPWR VPWR _04812_ sky130_fd_sc_hd__a22o_1
XFILLER_129_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_900 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09323_ net1109 net3884 net405 VGND VGND VPWR VPWR _01076_ sky130_fd_sc_hd__mux2_1
X_06535_ tag_array.tag1\[4\]\[6\] net1363 net1269 tag_array.tag1\[7\]\[6\] _03858_
+ VGND VGND VPWR VPWR _03859_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_138_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09254_ net764 net4167 net576 VGND VGND VPWR VPWR _01008_ sky130_fd_sc_hd__mux2_1
X_06466_ tag_array.tag1\[13\]\[0\] net1579 net1483 tag_array.tag1\[14\]\[0\] VGND
+ VGND VPWR VPWR _03796_ sky130_fd_sc_hd__a22o_1
XFILLER_139_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08205_ net778 net4206 net799 VGND VGND VPWR VPWR _00199_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09185_ net738 net3138 net628 VGND VGND VPWR VPWR _00939_ sky130_fd_sc_hd__mux2_1
X_06397_ tag_array.tag0\[12\]\[19\] net1405 net1311 tag_array.tag0\[15\]\[19\] _03732_
+ VGND VGND VPWR VPWR _03733_ sky130_fd_sc_hd__a221o_1
XFILLER_135_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_151_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08136_ data_array.data1\[5\]\[63\] net1553 net1457 data_array.data1\[6\]\[63\] VGND
+ VGND VPWR VPWR _05314_ sky130_fd_sc_hd__a22o_1
XFILLER_181_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_151_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08067_ _05250_ _05251_ VGND VGND VPWR VPWR _00115_ sky130_fd_sc_hd__or2_1
XFILLER_107_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_112_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_654 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07018_ data_array.data0\[5\]\[25\] net1519 net1423 data_array.data0\[6\]\[25\] VGND
+ VGND VPWR VPWR _04298_ sky130_fd_sc_hd__a22o_1
XFILLER_68_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2530 tag_array.tag0\[1\]\[5\] VGND VGND VPWR VPWR net4181 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2541 tag_array.tag0\[8\]\[6\] VGND VGND VPWR VPWR net4192 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2552 data_array.data0\[11\]\[27\] VGND VGND VPWR VPWR net4203 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2563 data_array.data0\[7\]\[25\] VGND VGND VPWR VPWR net4214 sky130_fd_sc_hd__dlygate4sd3_1
X_08969_ net888 net3059 net427 VGND VGND VPWR VPWR _00725_ sky130_fd_sc_hd__mux2_1
Xhold2574 data_array.data1\[14\]\[45\] VGND VGND VPWR VPWR net4225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1840 data_array.data1\[13\]\[21\] VGND VGND VPWR VPWR net3491 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_124_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2585 data_array.data0\[10\]\[33\] VGND VGND VPWR VPWR net4236 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1851 data_array.data0\[10\]\[61\] VGND VGND VPWR VPWR net3502 sky130_fd_sc_hd__dlygate4sd3_1
X_11980_ clknet_leaf_221_clk _00788_ VGND VGND VPWR VPWR data_array.data0\[4\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2596 tag_array.tag0\[13\]\[18\] VGND VGND VPWR VPWR net4247 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_151_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1862 tag_array.tag0\[6\]\[22\] VGND VGND VPWR VPWR net3513 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1873 data_array.data1\[7\]\[8\] VGND VGND VPWR VPWR net3524 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1884 tag_array.tag1\[11\]\[9\] VGND VGND VPWR VPWR net3535 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10931_ net1017 net4530 net528 VGND VGND VPWR VPWR _02676_ sky130_fd_sc_hd__mux2_1
Xhold1895 tag_array.tag0\[12\]\[18\] VGND VGND VPWR VPWR net3546 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_95_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_158_3407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13650_ clknet_leaf_119_clk _02279_ VGND VGND VPWR VPWR data_array.data1\[15\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10862_ net1038 net3520 net519 VGND VGND VPWR VPWR _02607_ sky130_fd_sc_hd__mux2_1
XFILLER_182_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_175_3721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_175_3732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12601_ clknet_leaf_144_clk _01295_ VGND VGND VPWR VPWR tag_array.tag0\[0\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_13581_ clknet_leaf_0_clk _02210_ VGND VGND VPWR VPWR data_array.data0\[9\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_25_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10793_ net1781 net1056 net505 VGND VGND VPWR VPWR _02538_ sky130_fd_sc_hd__mux2_1
XFILLER_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12532_ clknet_leaf_231_clk _01226_ VGND VGND VPWR VPWR tag_array.tag1\[11\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_158_938 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12463_ clknet_leaf_70_clk _01157_ VGND VGND VPWR VPWR data_array.data1\[9\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_172_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14202_ clknet_leaf_242_clk _02831_ VGND VGND VPWR VPWR data_array.data0\[2\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
X_11414_ clknet_leaf_48_clk _00224_ VGND VGND VPWR VPWR data_array.data0\[0\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_137_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12394_ clknet_leaf_94_clk _01088_ VGND VGND VPWR VPWR data_array.data0\[14\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_14133_ clknet_leaf_20_clk _02762_ VGND VGND VPWR VPWR data_array.data0\[1\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_137_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11345_ net915 net3804 net801 VGND VGND VPWR VPWR _03088_ sky130_fd_sc_hd__mux2_1
XFILLER_125_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14064_ clknet_leaf_123_clk _02693_ VGND VGND VPWR VPWR data_array.data1\[6\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
X_11276_ net925 net2379 net673 VGND VGND VPWR VPWR _03019_ sky130_fd_sc_hd__mux2_1
XFILLER_125_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13015_ clknet_leaf_70_clk _01709_ VGND VGND VPWR VPWR data_array.data0\[3\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_79_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10227_ net897 net3056 net354 VGND VGND VPWR VPWR _01974_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10158_ net913 net2809 net367 VGND VGND VPWR VPWR _01906_ sky130_fd_sc_hd__mux2_1
XFILLER_0_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_50_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_50_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10089_ net1880 net767 net638 VGND VGND VPWR VPWR _01838_ sky130_fd_sc_hd__mux2_1
X_13917_ clknet_leaf_229_clk _02546_ VGND VGND VPWR VPWR data_array.data1\[4\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13848_ clknet_leaf_214_clk _02477_ VGND VGND VPWR VPWR data_array.data1\[3\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13779_ clknet_leaf_36_clk _02408_ VGND VGND VPWR VPWR data_array.data1\[2\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_06320_ tag_array.tag0\[8\]\[12\] net1407 net1313 tag_array.tag0\[11\]\[12\] _03662_
+ VGND VGND VPWR VPWR _03663_ sky130_fd_sc_hd__a221o_1
XFILLER_128_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06251_ net1184 _03595_ _03599_ net1232 VGND VGND VPWR VPWR _03601_ sky130_fd_sc_hd__a22o_1
XFILLER_175_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_4_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_4_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_175_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06182_ tag_array.valid1\[5\] net1557 net1461 tag_array.valid1\[6\] VGND VGND VPWR
+ VPWR _03538_ sky130_fd_sc_hd__a22o_1
XFILLER_184_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold403 data_array.data1\[1\]\[32\] VGND VGND VPWR VPWR net2054 sky130_fd_sc_hd__dlygate4sd3_1
Xhold414 data_array.data0\[8\]\[35\] VGND VGND VPWR VPWR net2065 sky130_fd_sc_hd__dlygate4sd3_1
Xhold425 data_array.data0\[6\]\[9\] VGND VGND VPWR VPWR net2076 sky130_fd_sc_hd__dlygate4sd3_1
Xhold436 data_array.data0\[8\]\[44\] VGND VGND VPWR VPWR net2087 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold447 tag_array.tag0\[10\]\[9\] VGND VGND VPWR VPWR net2098 sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 data_array.data1\[8\]\[27\] VGND VGND VPWR VPWR net2109 sky130_fd_sc_hd__dlygate4sd3_1
X_09941_ net1064 net4510 net376 VGND VGND VPWR VPWR _01690_ sky130_fd_sc_hd__mux2_1
XFILLER_116_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold469 tag_array.tag0\[15\]\[23\] VGND VGND VPWR VPWR net2120 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout905 _05522_ VGND VGND VPWR VPWR net905 sky130_fd_sc_hd__buf_1
XFILLER_98_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout916 _05516_ VGND VGND VPWR VPWR net916 sky130_fd_sc_hd__clkbuf_2
Xfanout927 _05512_ VGND VGND VPWR VPWR net927 sky130_fd_sc_hd__buf_1
XFILLER_48_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09872_ net983 net4264 net378 VGND VGND VPWR VPWR _01622_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_70_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout938 net939 VGND VGND VPWR VPWR net938 sky130_fd_sc_hd__clkbuf_2
Xfanout949 _05500_ VGND VGND VPWR VPWR net949 sky130_fd_sc_hd__buf_1
XFILLER_38_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1103 data_array.data1\[6\]\[57\] VGND VGND VPWR VPWR net2754 sky130_fd_sc_hd__dlygate4sd3_1
X_08823_ net3589 net955 net449 VGND VGND VPWR VPWR _00581_ sky130_fd_sc_hd__mux2_1
Xhold1114 data_array.data0\[15\]\[25\] VGND VGND VPWR VPWR net2765 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1125 tag_array.tag0\[11\]\[0\] VGND VGND VPWR VPWR net2776 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1136 data_array.data1\[0\]\[22\] VGND VGND VPWR VPWR net2787 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1147 data_array.data1\[15\]\[0\] VGND VGND VPWR VPWR net2798 sky130_fd_sc_hd__dlygate4sd3_1
X_08754_ net707 net2629 net460 VGND VGND VPWR VPWR _00513_ sky130_fd_sc_hd__mux2_1
X_05966_ data_array.rdata0\[45\] net847 net1146 VGND VGND VPWR VPWR _03438_ sky130_fd_sc_hd__o21a_1
Xhold1158 data_array.data0\[11\]\[49\] VGND VGND VPWR VPWR net2809 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1169 data_array.data1\[0\]\[20\] VGND VGND VPWR VPWR net2820 sky130_fd_sc_hd__dlygate4sd3_1
X_07705_ data_array.data1\[13\]\[24\] net1586 net1490 data_array.data1\[14\]\[24\]
+ VGND VGND VPWR VPWR _04922_ sky130_fd_sc_hd__a22o_1
XFILLER_38_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08685_ net2482 net782 net486 VGND VGND VPWR VPWR _00444_ sky130_fd_sc_hd__mux2_1
X_05897_ data_array.rdata0\[22\] net847 net1143 VGND VGND VPWR VPWR _03392_ sky130_fd_sc_hd__o21a_1
XFILLER_53_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_92_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_92_clk sky130_fd_sc_hd__clkbuf_8
X_07636_ net1190 _04853_ _04857_ net1616 VGND VGND VPWR VPWR _04860_ sky130_fd_sc_hd__a22o_1
XFILLER_14_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_68_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07567_ data_array.data1\[12\]\[11\] net1384 net1290 data_array.data1\[15\]\[11\]
+ _04796_ VGND VGND VPWR VPWR _04797_ sky130_fd_sc_hd__a221o_1
X_09306_ net757 net4551 net551 VGND VGND VPWR VPWR _01060_ sky130_fd_sc_hd__mux2_1
XFILLER_179_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06518_ tag_array.tag1\[8\]\[5\] net1420 net1326 tag_array.tag1\[11\]\[5\] _03842_
+ VGND VGND VPWR VPWR _03843_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_153_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07498_ data_array.data1\[1\]\[5\] net1551 net1455 data_array.data1\[2\]\[5\] VGND
+ VGND VPWR VPWR _04734_ sky130_fd_sc_hd__a22o_1
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09237_ net733 net2312 net645 VGND VGND VPWR VPWR _00991_ sky130_fd_sc_hd__mux2_1
X_06449_ net1232 _03775_ _03779_ net1184 VGND VGND VPWR VPWR _03781_ sky130_fd_sc_hd__a22o_1
XFILLER_154_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09168_ net870 net3424 net576 VGND VGND VPWR VPWR _00922_ sky130_fd_sc_hd__mux2_1
XFILLER_5_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08119_ data_array.data1\[4\]\[61\] net1354 net1260 data_array.data1\[7\]\[61\] _05298_
+ VGND VGND VPWR VPWR _05299_ sky130_fd_sc_hd__a221o_1
XFILLER_162_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09099_ net888 net3510 net411 VGND VGND VPWR VPWR _00853_ sky130_fd_sc_hd__mux2_1
XFILLER_123_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11130_ net997 net3385 net544 VGND VGND VPWR VPWR _02873_ sky130_fd_sc_hd__mux2_1
XFILLER_122_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold970 tag_array.tag1\[11\]\[10\] VGND VGND VPWR VPWR net2621 sky130_fd_sc_hd__dlygate4sd3_1
Xhold981 data_array.data0\[2\]\[17\] VGND VGND VPWR VPWR net2632 sky130_fd_sc_hd__dlygate4sd3_1
X_11061_ net1953 net1018 net330 VGND VGND VPWR VPWR _02804_ sky130_fd_sc_hd__mux2_1
Xhold992 data_array.data0\[13\]\[10\] VGND VGND VPWR VPWR net2643 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_168_3591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10012_ net1038 net3120 net556 VGND VGND VPWR VPWR _01761_ sky130_fd_sc_hd__mux2_1
XFILLER_49_627 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2360 data_array.data1\[3\]\[46\] VGND VGND VPWR VPWR net4011 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_95_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2371 tag_array.tag0\[12\]\[4\] VGND VGND VPWR VPWR net4022 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2382 data_array.data0\[11\]\[41\] VGND VGND VPWR VPWR net4033 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_92_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2393 data_array.data0\[7\]\[29\] VGND VGND VPWR VPWR net4044 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1670 data_array.data1\[5\]\[48\] VGND VGND VPWR VPWR net3321 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_151_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1681 data_array.data0\[6\]\[17\] VGND VGND VPWR VPWR net3332 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_151_74 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11963_ clknet_leaf_217_clk _00771_ VGND VGND VPWR VPWR data_array.data0\[4\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1692 tag_array.tag1\[12\]\[1\] VGND VGND VPWR VPWR net3343 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_83_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_83_clk sky130_fd_sc_hd__clkbuf_8
X_13702_ clknet_leaf_121_clk _02331_ VGND VGND VPWR VPWR data_array.data1\[15\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
X_10914_ net1085 net2943 net526 VGND VGND VPWR VPWR _02659_ sky130_fd_sc_hd__mux2_1
X_11894_ clknet_leaf_264_clk _00702_ VGND VGND VPWR VPWR data_array.data0\[5\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13633_ clknet_leaf_207_clk _02262_ VGND VGND VPWR VPWR data_array.data0\[9\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
X_10845_ net1104 net4239 net514 VGND VGND VPWR VPWR _02590_ sky130_fd_sc_hd__mux2_1
XFILLER_60_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10776_ net870 net2439 net500 VGND VGND VPWR VPWR _02521_ sky130_fd_sc_hd__mux2_1
X_13564_ clknet_leaf_211_clk _02193_ VGND VGND VPWR VPWR data_array.data1\[0\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_157_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12515_ clknet_leaf_172_clk _01209_ VGND VGND VPWR VPWR lru_array.lru_mem\[10\] sky130_fd_sc_hd__dfxtp_1
X_13495_ clknet_leaf_31_clk _00130_ VGND VGND VPWR VPWR dirty_way1 sky130_fd_sc_hd__dfxtp_2
XFILLER_157_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12446_ clknet_leaf_175_clk _01140_ VGND VGND VPWR VPWR lru_array.lru_mem\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_126_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12377_ clknet_leaf_52_clk _00054_ VGND VGND VPWR VPWR data_array.rdata0\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_126_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11328_ net980 net4015 net795 VGND VGND VPWR VPWR _03071_ sky130_fd_sc_hd__mux2_1
X_14116_ clknet_leaf_29_clk _02745_ VGND VGND VPWR VPWR data_array.data0\[1\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_114_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14047_ clknet_leaf_204_clk _02676_ VGND VGND VPWR VPWR data_array.data1\[6\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_11259_ net994 net4596 net680 VGND VGND VPWR VPWR _03002_ sky130_fd_sc_hd__mux2_1
XFILLER_68_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05820_ _03258_ _03271_ _03272_ _03279_ VGND VGND VPWR VPWR _03337_ sky130_fd_sc_hd__or4_1
XFILLER_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_89_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_167_Right_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05751_ _03256_ _03257_ _03262_ _03267_ VGND VGND VPWR VPWR _03268_ sky130_fd_sc_hd__or4_1
XFILLER_35_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_74_clk clknet_5_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_74_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_35_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08470_ net1728 net665 VGND VGND VPWR VPWR _00286_ sky130_fd_sc_hd__or2_1
X_05682_ fsm.tag_out0\[5\] net4 VGND VGND VPWR VPWR _03199_ sky130_fd_sc_hd__and2b_1
XFILLER_35_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07421_ data_array.data0\[5\]\[62\] net1602 net1506 data_array.data0\[6\]\[62\] VGND
+ VGND VPWR VPWR _04664_ sky130_fd_sc_hd__a22o_1
XFILLER_63_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07352_ _04600_ _04601_ VGND VGND VPWR VPWR _00050_ sky130_fd_sc_hd__or2_1
XFILLER_148_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06303_ tag_array.tag0\[1\]\[10\] net1595 net1499 tag_array.tag0\[2\]\[10\] VGND
+ VGND VPWR VPWR _03648_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_100_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07283_ data_array.data0\[4\]\[49\] net1389 net1295 data_array.data0\[7\]\[49\] _04538_
+ VGND VGND VPWR VPWR _04539_ sky130_fd_sc_hd__a221o_1
X_09022_ net2200 net936 net423 VGND VGND VPWR VPWR _00777_ sky130_fd_sc_hd__mux2_1
XFILLER_136_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06234_ tag_array.tag0\[4\]\[4\] net1371 net1277 tag_array.tag0\[7\]\[4\] _03584_
+ VGND VGND VPWR VPWR _03585_ sky130_fd_sc_hd__a221o_1
XFILLER_148_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold200 data_array.data1\[0\]\[61\] VGND VGND VPWR VPWR net1851 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06165_ net28 net29 VGND VGND VPWR VPWR _03522_ sky130_fd_sc_hd__and2_1
Xhold211 data_array.data1\[1\]\[18\] VGND VGND VPWR VPWR net1862 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold222 data_array.data1\[1\]\[19\] VGND VGND VPWR VPWR net1873 sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 data_array.data0\[0\]\[48\] VGND VGND VPWR VPWR net1884 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 data_array.data0\[8\]\[48\] VGND VGND VPWR VPWR net1895 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold255 data_array.data0\[0\]\[12\] VGND VGND VPWR VPWR net1906 sky130_fd_sc_hd__dlygate4sd3_1
X_06096_ data_array.rdata0\[11\] net1140 net1114 data_array.rdata1\[11\] VGND VGND
+ VPWR VPWR net265 sky130_fd_sc_hd__a22o_1
XFILLER_171_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold266 data_array.data1\[4\]\[34\] VGND VGND VPWR VPWR net1917 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold277 data_array.data0\[1\]\[3\] VGND VGND VPWR VPWR net1928 sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 data_array.data0\[4\]\[16\] VGND VGND VPWR VPWR net1939 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout702 net703 VGND VGND VPWR VPWR net702 sky130_fd_sc_hd__clkbuf_2
X_09924_ net712 net4380 net602 VGND VGND VPWR VPWR _01674_ sky130_fd_sc_hd__mux2_1
XFILLER_131_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold299 data_array.data0\[8\]\[42\] VGND VGND VPWR VPWR net1950 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_59_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout713 _05405_ VGND VGND VPWR VPWR net713 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout724 _05399_ VGND VGND VPWR VPWR net724 sky130_fd_sc_hd__clkbuf_2
Xfanout735 net737 VGND VGND VPWR VPWR net735 sky130_fd_sc_hd__clkbuf_2
XFILLER_131_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout746 _05387_ VGND VGND VPWR VPWR net746 sky130_fd_sc_hd__clkbuf_2
X_09855_ net1049 net2854 net383 VGND VGND VPWR VPWR _01605_ sky130_fd_sc_hd__mux2_1
Xfanout757 _05383_ VGND VGND VPWR VPWR net757 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_146_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout768 net769 VGND VGND VPWR VPWR net768 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_146_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout779 net780 VGND VGND VPWR VPWR net779 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08806_ net1883 net1022 net443 VGND VGND VPWR VPWR _00564_ sky130_fd_sc_hd__mux2_1
X_06998_ net1197 _04273_ _04277_ net1623 VGND VGND VPWR VPWR _04280_ sky130_fd_sc_hd__a22o_1
X_09786_ net1064 net4432 net390 VGND VGND VPWR VPWR _01537_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Left_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05949_ data_array.rdata1\[39\] net828 net837 VGND VGND VPWR VPWR _03427_ sky130_fd_sc_hd__a21o_1
X_08737_ net775 net3225 net458 VGND VGND VPWR VPWR _00496_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_134_Right_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_65_clk clknet_5_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_65_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_124_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08668_ net750 net2537 net501 VGND VGND VPWR VPWR _00427_ sky130_fd_sc_hd__mux2_1
XFILLER_14_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07619_ data_array.data1\[5\]\[16\] net1545 net1449 data_array.data1\[6\]\[16\] VGND
+ VGND VPWR VPWR _04844_ sky130_fd_sc_hd__a22o_1
X_08599_ net729 net3948 net535 VGND VGND VPWR VPWR _00358_ sky130_fd_sc_hd__mux2_1
XFILLER_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10630_ net2209 net942 net473 VGND VGND VPWR VPWR _02375_ sky130_fd_sc_hd__mux2_1
XFILLER_14_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10561_ net960 net4514 net457 VGND VGND VPWR VPWR _02306_ sky130_fd_sc_hd__mux2_1
X_12300_ clknet_leaf_133_clk _01058_ VGND VGND VPWR VPWR tag_array.tag1\[12\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13280_ clknet_leaf_10_clk _01910_ VGND VGND VPWR VPWR data_array.data0\[11\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
X_10492_ net976 net3016 net349 VGND VGND VPWR VPWR _02237_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12231_ clknet_leaf_147_clk _00160_ VGND VGND VPWR VPWR fsm.tag_out1\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12162_ clknet_leaf_160_clk _00970_ VGND VGND VPWR VPWR tag_array.tag0\[13\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_943 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11113_ net1066 net2874 net548 VGND VGND VPWR VPWR _02856_ sky130_fd_sc_hd__mux2_1
XFILLER_146_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12093_ clknet_leaf_240_clk _00901_ VGND VGND VPWR VPWR data_array.data1\[14\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_49_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11044_ net2119 net1084 net328 VGND VGND VPWR VPWR _02787_ sky130_fd_sc_hd__mux2_1
XFILLER_118_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_183_3875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1025 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2190 data_array.data1\[7\]\[44\] VGND VGND VPWR VPWR net3841 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_101_Right_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_56_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_56_clk sky130_fd_sc_hd__clkbuf_8
X_12995_ clknet_leaf_112_clk _01689_ VGND VGND VPWR VPWR data_array.data0\[3\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_855 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11946_ clknet_leaf_127_clk _00754_ VGND VGND VPWR VPWR data_array.data0\[4\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_55_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11877_ clknet_leaf_63_clk _00685_ VGND VGND VPWR VPWR data_array.data0\[5\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_13616_ clknet_leaf_260_clk _02245_ VGND VGND VPWR VPWR data_array.data0\[9\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_45_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10828_ net2789 net918 net508 VGND VGND VPWR VPWR _02573_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13547_ clknet_leaf_83_clk _02176_ VGND VGND VPWR VPWR data_array.data1\[0\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_71_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10759_ net937 net3304 net496 VGND VGND VPWR VPWR _02504_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_41_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13478_ clknet_leaf_158_clk _02108_ VGND VGND VPWR VPWR tag_array.tag0\[15\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_145_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12429_ clknet_leaf_39_clk _01123_ VGND VGND VPWR VPWR data_array.data0\[14\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput305 net305 VGND VGND VPWR VPWR mem_wdata[48] sky130_fd_sc_hd__buf_2
Xoutput316 net316 VGND VGND VPWR VPWR mem_wdata[58] sky130_fd_sc_hd__buf_2
Xoutput327 net327 VGND VGND VPWR VPWR mem_write sky130_fd_sc_hd__buf_2
XFILLER_5_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07970_ data_array.data1\[8\]\[48\] net1397 net1303 data_array.data1\[11\]\[48\]
+ _05162_ VGND VGND VPWR VPWR _05163_ sky130_fd_sc_hd__a221o_1
X_06921_ net1624 _04203_ _04207_ net1195 VGND VGND VPWR VPWR _04210_ sky130_fd_sc_hd__a22o_1
XFILLER_171_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_1023 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09640_ net726 net2669 net617 VGND VGND VPWR VPWR _01392_ sky130_fd_sc_hd__mux2_1
X_06852_ data_array.data0\[12\]\[10\] net1411 net1317 data_array.data0\[15\]\[10\]
+ _04146_ VGND VGND VPWR VPWR _04147_ sky130_fd_sc_hd__a221o_1
X_05803_ _03316_ _03317_ _03318_ _03319_ VGND VGND VPWR VPWR _03320_ sky130_fd_sc_hd__or4_4
XFILLER_49_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09571_ net1064 net3881 net398 VGND VGND VPWR VPWR _01323_ sky130_fd_sc_hd__mux2_1
X_06783_ data_array.data0\[5\]\[4\] net1581 net1485 data_array.data0\[6\]\[4\] VGND
+ VGND VPWR VPWR _04084_ sky130_fd_sc_hd__a22o_1
XFILLER_83_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_47_clk clknet_5_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_47_clk sky130_fd_sc_hd__clkbuf_8
X_08522_ net821 net812 net854 _05352_ VGND VGND VPWR VPWR _05586_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_141_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05734_ net21 fsm.tag_out1\[21\] VGND VGND VPWR VPWR _03251_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_141_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08453_ net1866 net872 net692 VGND VGND VPWR VPWR _00280_ sky130_fd_sc_hd__mux2_1
XFILLER_51_633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05665_ fsm.tag_out0\[4\] net3 VGND VGND VPWR VPWR _03182_ sky130_fd_sc_hd__and2b_1
XFILLER_168_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07404_ data_array.data0\[0\]\[60\] net1411 net1317 data_array.data0\[3\]\[60\] _04648_
+ VGND VGND VPWR VPWR _04649_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_82_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08384_ net2053 net964 net693 VGND VGND VPWR VPWR _00257_ sky130_fd_sc_hd__mux2_1
X_07335_ data_array.data0\[13\]\[54\] net1547 net1451 data_array.data0\[14\]\[54\]
+ VGND VGND VPWR VPWR _04586_ sky130_fd_sc_hd__a22o_1
XFILLER_137_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07266_ data_array.data0\[8\]\[48\] net1391 net1297 data_array.data0\[11\]\[48\]
+ _04522_ VGND VGND VPWR VPWR _04523_ sky130_fd_sc_hd__a221o_1
X_09005_ net1868 net1006 net420 VGND VGND VPWR VPWR _00760_ sky130_fd_sc_hd__mux2_1
X_06217_ net1625 _03563_ _03567_ net1199 VGND VGND VPWR VPWR _03570_ sky130_fd_sc_hd__a22o_1
XFILLER_164_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07197_ net1167 _04455_ _04459_ net1215 VGND VGND VPWR VPWR _04461_ sky130_fd_sc_hd__a22o_1
XFILLER_118_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06148_ data_array.rdata0\[63\] net1137 net1118 data_array.rdata1\[63\] VGND VGND
+ VPWR VPWR net322 sky130_fd_sc_hd__a22o_1
XFILLER_133_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_148_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06079_ net1160 net22 fsm.tag_out1\[22\] net1131 VGND VGND VPWR VPWR _03503_ sky130_fd_sc_hd__a22o_1
Xfanout510 net511 VGND VGND VPWR VPWR net510 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1508 net1510 VGND VGND VPWR VPWR net1508 sky130_fd_sc_hd__clkbuf_4
Xfanout1519 net1521 VGND VGND VPWR VPWR net1519 sky130_fd_sc_hd__clkbuf_4
Xfanout521 net522 VGND VGND VPWR VPWR net521 sky130_fd_sc_hd__buf_2
X_09907_ net781 net3996 net602 VGND VGND VPWR VPWR _01657_ sky130_fd_sc_hd__mux2_1
XFILLER_99_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout532 net534 VGND VGND VPWR VPWR net532 sky130_fd_sc_hd__clkbuf_8
Xfanout543 net547 VGND VGND VPWR VPWR net543 sky130_fd_sc_hd__clkbuf_8
XFILLER_76_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout554 net560 VGND VGND VPWR VPWR net554 sky130_fd_sc_hd__buf_4
XFILLER_76_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout565 _05593_ VGND VGND VPWR VPWR net565 sky130_fd_sc_hd__buf_4
XFILLER_47_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout576 net577 VGND VGND VPWR VPWR net576 sky130_fd_sc_hd__buf_4
Xfanout587 net590 VGND VGND VPWR VPWR net587 sky130_fd_sc_hd__buf_2
X_09838_ net856 net3914 net388 VGND VGND VPWR VPWR _01589_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_161_3458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout598 _05586_ VGND VGND VPWR VPWR net598 sky130_fd_sc_hd__buf_2
XFILLER_46_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09769_ net2706 net711 net663 VGND VGND VPWR VPWR _01521_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_122_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_38_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_38_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_122_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ clknet_leaf_247_clk _00608_ VGND VGND VPWR VPWR data_array.data0\[7\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12780_ clknet_leaf_108_clk _01474_ VGND VGND VPWR VPWR tag_array.tag0\[6\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_162_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11731_ clknet_leaf_185_clk _00539_ VGND VGND VPWR VPWR tag_array.tag0\[9\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_942 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14450_ clknet_leaf_8_clk _03073_ VGND VGND VPWR VPWR data_array.data1\[7\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_25_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ clknet_leaf_192_clk _00470_ VGND VGND VPWR VPWR tag_array.tag1\[1\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13401_ clknet_leaf_228_clk _02031_ VGND VGND VPWR VPWR data_array.data1\[8\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_54_Left_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10613_ net2705 net1008 net466 VGND VGND VPWR VPWR _02358_ sky130_fd_sc_hd__mux2_1
X_14381_ clknet_leaf_39_clk _03004_ VGND VGND VPWR VPWR data_array.data1\[10\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_11593_ clknet_leaf_142_clk _00401_ VGND VGND VPWR VPWR tag_array.tag1\[4\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10544_ net1031 net3635 net463 VGND VGND VPWR VPWR _02289_ sky130_fd_sc_hd__mux2_1
X_13332_ clknet_leaf_260_clk _01962_ VGND VGND VPWR VPWR data_array.data0\[10\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_109_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13263_ clknet_leaf_114_clk _01893_ VGND VGND VPWR VPWR data_array.data0\[11\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
X_10475_ net1046 net2920 net346 VGND VGND VPWR VPWR _02220_ sky130_fd_sc_hd__mux2_1
XFILLER_142_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12214_ clknet_leaf_152_clk _00144_ VGND VGND VPWR VPWR fsm.tag_out0\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_155_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13194_ clknet_leaf_49_clk _00088_ VGND VGND VPWR VPWR data_array.rdata1\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_151_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12145_ clknet_leaf_170_clk _00953_ VGND VGND VPWR VPWR tag_array.tag0\[13\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_151_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_63_Left_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12076_ clknet_leaf_24_clk _00884_ VGND VGND VPWR VPWR data_array.data1\[14\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_89_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11027_ net2404 net895 net338 VGND VGND VPWR VPWR _02771_ sky130_fd_sc_hd__mux2_1
XFILLER_49_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_86_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_29_clk clknet_5_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_64_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12978_ clknet_leaf_153_clk _01672_ VGND VGND VPWR VPWR tag_array.tag0\[4\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11929_ clknet_leaf_48_clk _00737_ VGND VGND VPWR VPWR data_array.data0\[4\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_43_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_72_Left_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_17 _03477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_28 _05417_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_39 net472 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07120_ net1168 _04385_ _04389_ net1216 VGND VGND VPWR VPWR _04391_ sky130_fd_sc_hd__a22o_1
XFILLER_174_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07051_ data_array.data0\[1\]\[28\] net1540 net1444 data_array.data0\[2\]\[28\] VGND
+ VGND VPWR VPWR _04328_ sky130_fd_sc_hd__a22o_1
XFILLER_161_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06002_ data_array.rdata0\[57\] net848 net1144 VGND VGND VPWR VPWR _03462_ sky130_fd_sc_hd__o21a_1
XFILLER_12_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput168 net168 VGND VGND VPWR VPWR cpu_rdata[12] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_58_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_81_Left_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput179 net179 VGND VGND VPWR VPWR cpu_rdata[22] sky130_fd_sc_hd__buf_2
XFILLER_142_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2904 data_array.data1\[7\]\[26\] VGND VGND VPWR VPWR net4555 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2915 tag_array.tag1\[14\]\[3\] VGND VGND VPWR VPWR net4566 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2926 data_array.data0\[15\]\[1\] VGND VGND VPWR VPWR net4577 sky130_fd_sc_hd__dlygate4sd3_1
X_07953_ data_array.data1\[1\]\[46\] net1524 net1428 data_array.data1\[2\]\[46\] VGND
+ VGND VPWR VPWR _05148_ sky130_fd_sc_hd__a22o_1
Xhold2937 data_array.data0\[6\]\[46\] VGND VGND VPWR VPWR net4588 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_101_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2948 data_array.data0\[10\]\[38\] VGND VGND VPWR VPWR net4599 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_143_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2959 tag_array.tag0\[7\]\[7\] VGND VGND VPWR VPWR net4610 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_143_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06904_ data_array.data0\[5\]\[15\] net1580 net1484 data_array.data0\[6\]\[15\] VGND
+ VGND VPWR VPWR _04194_ sky130_fd_sc_hd__a22o_1
X_07884_ data_array.data1\[4\]\[40\] net1415 net1321 data_array.data1\[7\]\[40\] _05084_
+ VGND VGND VPWR VPWR _05085_ sky130_fd_sc_hd__a221o_1
XFILLER_95_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09623_ net856 net3740 net396 VGND VGND VPWR VPWR _01375_ sky130_fd_sc_hd__mux2_1
XFILLER_110_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06835_ _04130_ _04131_ VGND VGND VPWR VPWR _00062_ sky130_fd_sc_hd__or2_1
XFILLER_95_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06766_ data_array.data0\[0\]\[2\] net1338 net1244 data_array.data0\[3\]\[2\] _04068_
+ VGND VGND VPWR VPWR _04069_ sky130_fd_sc_hd__a221o_1
X_09554_ net713 net4544 net618 VGND VGND VPWR VPWR _01307_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_90_Left_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08505_ net1714 net614 VGND VGND VPWR VPWR _00297_ sky130_fd_sc_hd__nand2b_1
X_05717_ _03135_ fsm.tag_out0\[1\] _03169_ _03170_ _03185_ VGND VGND VPWR VPWR _03234_
+ sky130_fd_sc_hd__a2111o_1
X_09485_ net789 net3407 net624 VGND VGND VPWR VPWR _01238_ sky130_fd_sc_hd__mux2_1
X_06697_ tag_array.tag1\[13\]\[21\] net1595 net1499 tag_array.tag1\[14\]\[21\] VGND
+ VGND VPWR VPWR _04006_ sky130_fd_sc_hd__a22o_1
XFILLER_23_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08436_ net148 net83 net1643 VGND VGND VPWR VPWR _05527_ sky130_fd_sc_hd__mux2_1
X_05648_ net32 fsm.tag_out0\[2\] VGND VGND VPWR VPWR _03165_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_22_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08367_ net123 net58 net1640 VGND VGND VPWR VPWR _05481_ sky130_fd_sc_hd__mux2_1
XFILLER_134_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07318_ net1170 _04565_ _04569_ net1218 VGND VGND VPWR VPWR _04571_ sky130_fd_sc_hd__a22o_1
X_08298_ net161 net96 net1638 VGND VGND VPWR VPWR _05435_ sky130_fd_sc_hd__mux2_1
X_07249_ data_array.data0\[1\]\[46\] net1532 net1436 data_array.data0\[2\]\[46\] VGND
+ VGND VPWR VPWR _04508_ sky130_fd_sc_hd__a22o_1
XFILLER_152_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_847 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10260_ net705 net3360 net598 VGND VGND VPWR VPWR _02007_ sky130_fd_sc_hd__mux2_1
XFILLER_124_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10191_ net1043 net3875 net354 VGND VGND VPWR VPWR _01938_ sky130_fd_sc_hd__mux2_1
Xfanout1305 net1306 VGND VGND VPWR VPWR net1305 sky130_fd_sc_hd__clkbuf_4
Xfanout1316 net1328 VGND VGND VPWR VPWR net1316 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_180_3812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1327 net1328 VGND VGND VPWR VPWR net1327 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_180_3823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1338 net1339 VGND VGND VPWR VPWR net1338 sky130_fd_sc_hd__clkbuf_4
Xfanout340 _03132_ VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__clkbuf_4
Xfanout351 _03131_ VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__buf_4
Xfanout1349 net1351 VGND VGND VPWR VPWR net1349 sky130_fd_sc_hd__clkbuf_4
Xfanout362 net363 VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__buf_4
X_13950_ clknet_leaf_215_clk _02579_ VGND VGND VPWR VPWR data_array.data1\[4\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout373 net374 VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__clkbuf_4
Xfanout384 net385 VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__clkbuf_8
XFILLER_59_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout395 net401 VGND VGND VPWR VPWR net395 sky130_fd_sc_hd__buf_4
X_12901_ clknet_leaf_205_clk _01595_ VGND VGND VPWR VPWR data_array.data0\[13\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_13881_ clknet_leaf_55_clk _02510_ VGND VGND VPWR VPWR data_array.data1\[3\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
X_12832_ clknet_leaf_227_clk _01526_ VGND VGND VPWR VPWR data_array.data0\[12\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_98_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12763_ clknet_leaf_179_clk _01457_ VGND VGND VPWR VPWR tag_array.tag0\[6\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_178_3774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_3785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ clknet_leaf_138_clk _00522_ VGND VGND VPWR VPWR tag_array.tag0\[9\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12694_ clknet_leaf_153_clk _01388_ VGND VGND VPWR VPWR tag_array.tag0\[8\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_14433_ clknet_leaf_253_clk _03056_ VGND VGND VPWR VPWR data_array.data1\[7\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11645_ clknet_leaf_33_clk _00453_ VGND VGND VPWR VPWR tag_array.tag1\[2\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_161_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput15 cpu_addr[22] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_2
X_14364_ clknet_leaf_42_clk _02987_ VGND VGND VPWR VPWR data_array.data1\[10\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11576_ clknet_leaf_128_clk _00384_ VGND VGND VPWR VPWR tag_array.tag1\[5\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput26 cpu_addr[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_4
XFILLER_122_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput37 cpu_wdata[12] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_1
Xinput48 cpu_wdata[22] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_1
XFILLER_128_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput59 cpu_wdata[32] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_1
X_13315_ clknet_leaf_92_clk _01945_ VGND VGND VPWR VPWR data_array.data0\[10\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_10527_ net1098 net4494 net455 VGND VGND VPWR VPWR _02272_ sky130_fd_sc_hd__mux2_1
XFILLER_143_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14295_ clknet_leaf_70_clk _02924_ VGND VGND VPWR VPWR data_array.data1\[11\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_182_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13246_ clknet_leaf_60_clk _01876_ VGND VGND VPWR VPWR data_array.data0\[11\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_10458_ _05415_ _05590_ VGND VGND VPWR VPWR _03131_ sky130_fd_sc_hd__nand2_1
XFILLER_170_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10389_ net2012 net1098 net667 VGND VGND VPWR VPWR _02135_ sky130_fd_sc_hd__mux2_1
X_13177_ clknet_leaf_49_clk _00069_ VGND VGND VPWR VPWR data_array.rdata1\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_112_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12128_ clknet_leaf_108_clk _00936_ VGND VGND VPWR VPWR tag_array.tag0\[12\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_36_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12059_ clknet_leaf_197_clk _00867_ VGND VGND VPWR VPWR data_array.data1\[14\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_38_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06620_ tag_array.tag1\[13\]\[14\] net1558 net1462 tag_array.tag1\[14\]\[14\] VGND
+ VGND VPWR VPWR _03936_ sky130_fd_sc_hd__a22o_1
XFILLER_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06551_ tag_array.tag1\[8\]\[8\] net1417 net1323 tag_array.tag1\[11\]\[8\] _03872_
+ VGND VGND VPWR VPWR _03873_ sky130_fd_sc_hd__a221o_1
XFILLER_33_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09270_ net701 net3863 net577 VGND VGND VPWR VPWR _01024_ sky130_fd_sc_hd__mux2_1
X_06482_ net1181 _03805_ _03809_ net1229 VGND VGND VPWR VPWR _03811_ sky130_fd_sc_hd__a22o_1
XFILLER_61_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08221_ net1650 net1162 net8 VGND VGND VPWR VPWR _05382_ sky130_fd_sc_hd__and3_1
XFILLER_166_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08152_ tag_array.dirty1\[4\] net1350 net1256 tag_array.dirty1\[7\] _05328_ VGND
+ VGND VPWR VPWR _05329_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_99_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07103_ data_array.data0\[0\]\[33\] net1396 net1302 data_array.data0\[3\]\[33\] _04374_
+ VGND VGND VPWR VPWR _04375_ sky130_fd_sc_hd__a221o_1
X_08083_ data_array.data1\[13\]\[58\] net1550 net1454 data_array.data1\[14\]\[58\]
+ VGND VGND VPWR VPWR _05266_ sky130_fd_sc_hd__a22o_1
Xclkload220 clknet_leaf_154_clk VGND VGND VPWR VPWR clkload220/Y sky130_fd_sc_hd__inv_6
Xclkload231 clknet_leaf_129_clk VGND VGND VPWR VPWR clkload231/Y sky130_fd_sc_hd__inv_6
Xclkbuf_leaf_9_clk clknet_5_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_8
Xclkload242 clknet_leaf_139_clk VGND VGND VPWR VPWR clkload242/Y sky130_fd_sc_hd__inv_8
Xclkbuf_5_15__f_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_5_15__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_07034_ data_array.data0\[9\]\[27\] net1555 net1459 data_array.data0\[10\]\[27\]
+ VGND VGND VPWR VPWR _04312_ sky130_fd_sc_hd__a22o_1
XFILLER_161_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2701 data_array.data1\[9\]\[40\] VGND VGND VPWR VPWR net4352 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2712 data_array.data0\[5\]\[27\] VGND VGND VPWR VPWR net4363 sky130_fd_sc_hd__dlygate4sd3_1
X_08985_ net1912 net1084 net418 VGND VGND VPWR VPWR _00740_ sky130_fd_sc_hd__mux2_1
Xhold2723 data_array.data1\[14\]\[57\] VGND VGND VPWR VPWR net4374 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_110_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2734 tag_array.tag0\[9\]\[19\] VGND VGND VPWR VPWR net4385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2745 data_array.data0\[13\]\[59\] VGND VGND VPWR VPWR net4396 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2756 data_array.data0\[13\]\[46\] VGND VGND VPWR VPWR net4407 sky130_fd_sc_hd__dlygate4sd3_1
X_07936_ data_array.data1\[13\]\[45\] net1540 net1444 data_array.data1\[14\]\[45\]
+ VGND VGND VPWR VPWR _05132_ sky130_fd_sc_hd__a22o_1
XFILLER_180_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2767 tag_array.tag1\[10\]\[15\] VGND VGND VPWR VPWR net4418 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2778 data_array.data0\[11\]\[4\] VGND VGND VPWR VPWR net4429 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_980 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2789 data_array.data1\[10\]\[24\] VGND VGND VPWR VPWR net4440 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07867_ net1631 _05063_ _05067_ net1205 VGND VGND VPWR VPWR _05070_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_119_Left_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09606_ net926 net4546 net394 VGND VGND VPWR VPWR _01358_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06818_ data_array.data0\[13\]\[7\] net1601 net1505 data_array.data0\[14\]\[7\] VGND
+ VGND VPWR VPWR _04116_ sky130_fd_sc_hd__a22o_1
X_07798_ data_array.data1\[8\]\[32\] net1330 net1236 data_array.data1\[11\]\[32\]
+ _05006_ VGND VGND VPWR VPWR _05007_ sky130_fd_sc_hd__a221o_1
XFILLER_25_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09537_ net779 net3894 net618 VGND VGND VPWR VPWR _01290_ sky130_fd_sc_hd__mux2_1
X_06749_ data_array.data0\[12\]\[1\] net1333 net1239 data_array.data0\[15\]\[1\] _04052_
+ VGND VGND VPWR VPWR _04053_ sky130_fd_sc_hd__a221o_1
XFILLER_19_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09468_ net757 net3535 net658 VGND VGND VPWR VPWR _01221_ sky130_fd_sc_hd__mux2_1
XFILLER_25_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_156_3357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08419_ net1127 _05515_ VGND VGND VPWR VPWR _05516_ sky130_fd_sc_hd__and2_2
XFILLER_145_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09399_ net1070 net3931 net588 VGND VGND VPWR VPWR _01152_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_173_3682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11430_ clknet_leaf_59_clk _00240_ VGND VGND VPWR VPWR data_array.data0\[0\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_117_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_128_Left_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11361_ net1646 net3060 net539 VGND VGND VPWR VPWR _03104_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_134_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13100_ clknet_leaf_4_clk _01794_ VGND VGND VPWR VPWR data_array.data1\[13\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_98_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10312_ net1937 net914 net639 VGND VGND VPWR VPWR _02059_ sky130_fd_sc_hd__mux2_1
X_11292_ net863 net4097 net683 VGND VGND VPWR VPWR _03035_ sky130_fd_sc_hd__mux2_1
XFILLER_164_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14080_ clknet_leaf_13_clk _02709_ VGND VGND VPWR VPWR data_array.data1\[6\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_138_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13031_ clknet_leaf_23_clk _01725_ VGND VGND VPWR VPWR data_array.data0\[3\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
X_10243_ net770 net3083 net596 VGND VGND VPWR VPWR _01990_ sky130_fd_sc_hd__mux2_1
XFILLER_79_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1102 net1103 VGND VGND VPWR VPWR net1102 sky130_fd_sc_hd__clkbuf_2
X_10174_ net1109 net4246 net356 VGND VGND VPWR VPWR _01921_ sky130_fd_sc_hd__mux2_1
XFILLER_152_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1113 net1116 VGND VGND VPWR VPWR net1113 sky130_fd_sc_hd__buf_4
XFILLER_120_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1124 net1130 VGND VGND VPWR VPWR net1124 sky130_fd_sc_hd__buf_4
XFILLER_121_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1135 net1138 VGND VGND VPWR VPWR net1135 sky130_fd_sc_hd__buf_4
XFILLER_94_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1146 _03154_ VGND VGND VPWR VPWR net1146 sky130_fd_sc_hd__clkbuf_8
Xfanout1157 _03153_ VGND VGND VPWR VPWR net1157 sky130_fd_sc_hd__clkbuf_8
Xfanout1168 net1169 VGND VGND VPWR VPWR net1168 sky130_fd_sc_hd__buf_4
XFILLER_120_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1179 net1180 VGND VGND VPWR VPWR net1179 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_137_Left_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13933_ clknet_leaf_214_clk _02562_ VGND VGND VPWR VPWR data_array.data1\[4\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13864_ clknet_leaf_257_clk _02493_ VGND VGND VPWR VPWR data_array.data1\[3\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12815_ clknet_leaf_138_clk _01509_ VGND VGND VPWR VPWR tag_array.tag1\[0\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_13795_ clknet_leaf_248_clk _02424_ VGND VGND VPWR VPWR data_array.data1\[2\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_12746_ clknet_leaf_169_clk _01440_ VGND VGND VPWR VPWR tag_array.tag0\[5\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_176_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12677_ clknet_leaf_51_clk _01371_ VGND VGND VPWR VPWR data_array.data0\[15\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_13_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_146_Left_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14416_ clknet_leaf_227_clk _03039_ VGND VGND VPWR VPWR data_array.data1\[7\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_11628_ clknet_leaf_100_clk _00436_ VGND VGND VPWR VPWR tag_array.tag1\[3\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14347_ clknet_leaf_184_clk _00184_ _00192_ VGND VGND VPWR VPWR fsm.state\[3\] sky130_fd_sc_hd__dfrtp_1
X_11559_ clknet_leaf_97_clk _00367_ VGND VGND VPWR VPWR tag_array.tag1\[5\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_128_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold607 data_array.data0\[14\]\[10\] VGND VGND VPWR VPWR net2258 sky130_fd_sc_hd__dlygate4sd3_1
Xhold618 data_array.data0\[4\]\[62\] VGND VGND VPWR VPWR net2269 sky130_fd_sc_hd__dlygate4sd3_1
Xhold629 tag_array.tag0\[1\]\[21\] VGND VGND VPWR VPWR net2280 sky130_fd_sc_hd__dlygate4sd3_1
X_14278_ clknet_leaf_121_clk _02907_ VGND VGND VPWR VPWR data_array.data1\[12\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_38_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13229_ clknet_leaf_248_clk _01859_ VGND VGND VPWR VPWR data_array.data0\[11\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_40_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_560 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2008 data_array.data0\[13\]\[18\] VGND VGND VPWR VPWR net3659 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2019 tag_array.tag0\[5\]\[1\] VGND VGND VPWR VPWR net3670 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_155_Left_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_260_clk clknet_5_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_260_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold1307 data_array.data0\[14\]\[26\] VGND VGND VPWR VPWR net2958 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1318 data_array.data1\[3\]\[62\] VGND VGND VPWR VPWR net2969 sky130_fd_sc_hd__dlygate4sd3_1
X_05982_ data_array.rdata1\[50\] net828 net838 VGND VGND VPWR VPWR _03449_ sky130_fd_sc_hd__a21o_1
X_08770_ net745 net3514 net450 VGND VGND VPWR VPWR _00529_ sky130_fd_sc_hd__mux2_1
Xhold1329 data_array.data1\[2\]\[14\] VGND VGND VPWR VPWR net2980 sky130_fd_sc_hd__dlygate4sd3_1
X_07721_ data_array.data1\[8\]\[25\] net1330 net1236 data_array.data1\[11\]\[25\]
+ _04936_ VGND VGND VPWR VPWR _04937_ sky130_fd_sc_hd__a221o_1
XFILLER_38_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07652_ data_array.data1\[5\]\[19\] net1584 net1488 data_array.data1\[6\]\[19\] VGND
+ VGND VPWR VPWR _04874_ sky130_fd_sc_hd__a22o_1
XFILLER_81_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06603_ net1181 _03915_ _03919_ net1229 VGND VGND VPWR VPWR _03921_ sky130_fd_sc_hd__a22o_1
X_07583_ _04810_ _04811_ VGND VGND VPWR VPWR _00067_ sky130_fd_sc_hd__or2_1
XFILLER_179_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06534_ tag_array.tag1\[5\]\[6\] net1552 net1456 tag_array.tag1\[6\]\[6\] VGND VGND
+ VPWR VPWR _03858_ sky130_fd_sc_hd__a22o_1
X_09322_ _05414_ _05552_ VGND VGND VPWR VPWR _03123_ sky130_fd_sc_hd__or2_1
XFILLER_178_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09253_ net767 net2636 net571 VGND VGND VPWR VPWR _01007_ sky130_fd_sc_hd__mux2_1
X_06465_ tag_array.tag1\[0\]\[0\] net1385 net1291 tag_array.tag1\[3\]\[0\] _03794_
+ VGND VGND VPWR VPWR _03795_ sky130_fd_sc_hd__a221o_1
XFILLER_138_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08204_ fsm.tag_out1\[3\] net816 net808 fsm.tag_out0\[3\] _05370_ VGND VGND VPWR
+ VPWR _05371_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_79_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09184_ net744 net2778 net627 VGND VGND VPWR VPWR _00938_ sky130_fd_sc_hd__mux2_1
XFILLER_18_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06396_ tag_array.tag0\[13\]\[19\] net1613 net1517 tag_array.tag0\[14\]\[19\] VGND
+ VGND VPWR VPWR _03732_ sky130_fd_sc_hd__a22o_1
XFILLER_147_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08135_ data_array.data1\[12\]\[63\] net1361 net1267 data_array.data1\[15\]\[63\]
+ _05312_ VGND VGND VPWR VPWR _05313_ sky130_fd_sc_hd__a221o_1
XFILLER_174_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_151_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_1023 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_151_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08066_ net1168 _05245_ _05249_ net1216 VGND VGND VPWR VPWR _05251_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_112_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07017_ data_array.data0\[8\]\[25\] net1332 net1238 data_array.data0\[11\]\[25\]
+ _04296_ VGND VGND VPWR VPWR _04297_ sky130_fd_sc_hd__a221o_1
XFILLER_1_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2520 data_array.data1\[11\]\[19\] VGND VGND VPWR VPWR net4171 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_251_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_251_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold2531 tag_array.tag0\[3\]\[20\] VGND VGND VPWR VPWR net4182 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2542 data_array.data0\[10\]\[32\] VGND VGND VPWR VPWR net4193 sky130_fd_sc_hd__dlygate4sd3_1
X_08968_ net895 net4607 net428 VGND VGND VPWR VPWR _00724_ sky130_fd_sc_hd__mux2_1
XFILLER_25_1051 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2553 tag_array.tag1\[11\]\[12\] VGND VGND VPWR VPWR net4204 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2564 tag_array.tag1\[8\]\[20\] VGND VGND VPWR VPWR net4215 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1830 lru_array.lru_mem\[15\] VGND VGND VPWR VPWR net3481 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2575 data_array.data0\[7\]\[18\] VGND VGND VPWR VPWR net4226 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1841 data_array.data0\[12\]\[4\] VGND VGND VPWR VPWR net3492 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2586 tag_array.tag1\[6\]\[8\] VGND VGND VPWR VPWR net4237 sky130_fd_sc_hd__dlygate4sd3_1
X_07919_ data_array.data1\[12\]\[43\] net1378 net1284 data_array.data1\[15\]\[43\]
+ _05116_ VGND VGND VPWR VPWR _05117_ sky130_fd_sc_hd__a221o_1
Xhold1852 data_array.data1\[15\]\[26\] VGND VGND VPWR VPWR net3503 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2597 data_array.data1\[14\]\[59\] VGND VGND VPWR VPWR net4248 sky130_fd_sc_hd__dlygate4sd3_1
X_08899_ net909 net4562 net435 VGND VGND VPWR VPWR _00656_ sky130_fd_sc_hd__mux2_1
XFILLER_84_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1863 tag_array.tag0\[9\]\[12\] VGND VGND VPWR VPWR net3514 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1874 tag_array.dirty0\[5\] VGND VGND VPWR VPWR net3525 sky130_fd_sc_hd__dlygate4sd3_1
X_10930_ net1022 net3793 net527 VGND VGND VPWR VPWR _02675_ sky130_fd_sc_hd__mux2_1
XFILLER_95_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1885 tag_array.tag0\[11\]\[11\] VGND VGND VPWR VPWR net3536 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1896 tag_array.tag1\[11\]\[15\] VGND VGND VPWR VPWR net3547 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_158_3408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10861_ net1040 net2340 net514 VGND VGND VPWR VPWR _02606_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_175_3722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12600_ clknet_leaf_142_clk _01294_ VGND VGND VPWR VPWR tag_array.tag0\[0\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13580_ clknet_leaf_205_clk _02209_ VGND VGND VPWR VPWR data_array.data0\[9\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_10792_ net2116 net1062 net508 VGND VGND VPWR VPWR _02537_ sky130_fd_sc_hd__mux2_1
X_12531_ clknet_leaf_134_clk _01225_ VGND VGND VPWR VPWR tag_array.tag1\[11\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12462_ clknet_leaf_42_clk _01156_ VGND VGND VPWR VPWR data_array.data1\[9\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_14201_ clknet_leaf_52_clk _02830_ VGND VGND VPWR VPWR data_array.data0\[2\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
X_11413_ clknet_leaf_247_clk _00223_ VGND VGND VPWR VPWR data_array.data0\[0\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12393_ clknet_leaf_45_clk _01087_ VGND VGND VPWR VPWR data_array.data0\[14\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_153_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14132_ clknet_leaf_87_clk _02761_ VGND VGND VPWR VPWR data_array.data0\[1\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_181_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11344_ net918 net4336 net801 VGND VGND VPWR VPWR _03087_ sky130_fd_sc_hd__mux2_1
XFILLER_137_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14063_ clknet_leaf_238_clk _02692_ VGND VGND VPWR VPWR data_array.data1\[6\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
X_11275_ net931 net3190 net675 VGND VGND VPWR VPWR _03018_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_148_Right_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13014_ clknet_leaf_53_clk _01708_ VGND VGND VPWR VPWR data_array.data0\[3\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_10226_ net902 net2341 net356 VGND VGND VPWR VPWR _01973_ sky130_fd_sc_hd__mux2_1
XFILLER_3_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_242_clk clknet_5_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_242_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10157_ net917 net2495 net367 VGND VGND VPWR VPWR _01905_ sky130_fd_sc_hd__mux2_1
XFILLER_79_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_50_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10088_ net2913 net772 net642 VGND VGND VPWR VPWR _01837_ sky130_fd_sc_hd__mux2_1
XFILLER_94_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13916_ clknet_leaf_130_clk _02545_ VGND VGND VPWR VPWR data_array.data1\[4\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13847_ clknet_leaf_66_clk _02476_ VGND VGND VPWR VPWR data_array.data1\[3\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_18_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13778_ clknet_leaf_117_clk _02407_ VGND VGND VPWR VPWR data_array.data1\[2\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12729_ clknet_leaf_181_clk _01423_ VGND VGND VPWR VPWR tag_array.tag0\[7\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_148_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06250_ net1208 _03593_ _03597_ net1634 VGND VGND VPWR VPWR _03600_ sky130_fd_sc_hd__a22o_1
XFILLER_176_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06181_ tag_array.valid1\[8\] net1369 net1275 tag_array.valid1\[11\] _03536_ VGND
+ VGND VPWR VPWR _03537_ sky130_fd_sc_hd__a221o_1
Xhold404 tag_array.tag1\[1\]\[2\] VGND VGND VPWR VPWR net2055 sky130_fd_sc_hd__dlygate4sd3_1
Xhold415 data_array.data1\[8\]\[13\] VGND VGND VPWR VPWR net2066 sky130_fd_sc_hd__dlygate4sd3_1
Xhold426 data_array.data1\[1\]\[58\] VGND VGND VPWR VPWR net2077 sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 data_array.data1\[2\]\[18\] VGND VGND VPWR VPWR net2088 sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 tag_array.tag0\[13\]\[7\] VGND VGND VPWR VPWR net2099 sky130_fd_sc_hd__dlygate4sd3_1
Xhold459 data_array.data1\[1\]\[43\] VGND VGND VPWR VPWR net2110 sky130_fd_sc_hd__dlygate4sd3_1
X_09940_ net1068 net2411 net377 VGND VGND VPWR VPWR _01689_ sky130_fd_sc_hd__mux2_1
XFILLER_144_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout906 _05522_ VGND VGND VPWR VPWR net906 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_115_Right_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09871_ net987 net3161 net382 VGND VGND VPWR VPWR _01621_ sky130_fd_sc_hd__mux2_1
Xfanout917 _05516_ VGND VGND VPWR VPWR net917 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_70_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout928 net929 VGND VGND VPWR VPWR net928 sky130_fd_sc_hd__clkbuf_2
Xfanout939 _05506_ VGND VGND VPWR VPWR net939 sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_233_clk clknet_5_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_233_clk
+ sky130_fd_sc_hd__clkbuf_8
X_08822_ net2699 net957 net446 VGND VGND VPWR VPWR _00580_ sky130_fd_sc_hd__mux2_1
XFILLER_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1104 data_array.data0\[15\]\[53\] VGND VGND VPWR VPWR net2755 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1115 data_array.data0\[5\]\[50\] VGND VGND VPWR VPWR net2766 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1126 data_array.data1\[13\]\[61\] VGND VGND VPWR VPWR net2777 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1137 data_array.data0\[5\]\[30\] VGND VGND VPWR VPWR net2788 sky130_fd_sc_hd__dlygate4sd3_1
X_08753_ net710 net3893 net456 VGND VGND VPWR VPWR _00512_ sky130_fd_sc_hd__mux2_1
X_05965_ net137 net1156 _03436_ _03437_ VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__a22o_1
Xhold1148 data_array.data1\[6\]\[36\] VGND VGND VPWR VPWR net2799 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1159 data_array.data0\[14\]\[61\] VGND VGND VPWR VPWR net2810 sky130_fd_sc_hd__dlygate4sd3_1
X_07704_ _04920_ _04921_ VGND VGND VPWR VPWR _00079_ sky130_fd_sc_hd__or2_1
XFILLER_94_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05896_ net112 net1152 _03390_ _03391_ VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__a22o_1
XFILLER_53_300 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08684_ net1867 net786 net483 VGND VGND VPWR VPWR _00443_ sky130_fd_sc_hd__mux2_1
XFILLER_38_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07635_ data_array.data1\[4\]\[17\] net1336 net1242 data_array.data1\[7\]\[17\] _04858_
+ VGND VGND VPWR VPWR _04859_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_105_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07566_ data_array.data1\[13\]\[11\] net1574 net1478 data_array.data1\[14\]\[11\]
+ VGND VGND VPWR VPWR _04796_ sky130_fd_sc_hd__a22o_1
XFILLER_110_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09305_ net760 net2885 net552 VGND VGND VPWR VPWR _01059_ sky130_fd_sc_hd__mux2_1
X_06517_ tag_array.tag1\[9\]\[5\] net1611 net1515 tag_array.tag1\[10\]\[5\] VGND VGND
+ VPWR VPWR _03842_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_153_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07497_ data_array.data1\[8\]\[5\] net1360 net1266 data_array.data1\[11\]\[5\] _04732_
+ VGND VGND VPWR VPWR _04733_ sky130_fd_sc_hd__a221o_1
XFILLER_10_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09236_ net736 net2578 net645 VGND VGND VPWR VPWR _00990_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_170_3630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06448_ net1634 _03773_ _03777_ net1208 VGND VGND VPWR VPWR _03780_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09167_ net874 net4248 net573 VGND VGND VPWR VPWR _00921_ sky130_fd_sc_hd__mux2_1
X_06379_ tag_array.tag0\[8\]\[17\] net1405 net1311 tag_array.tag0\[11\]\[17\] _03716_
+ VGND VGND VPWR VPWR _03717_ sky130_fd_sc_hd__a221o_1
XFILLER_163_931 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08118_ data_array.data1\[5\]\[61\] net1545 net1449 data_array.data1\[6\]\[61\] VGND
+ VGND VPWR VPWR _05298_ sky130_fd_sc_hd__a22o_1
XFILLER_79_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09098_ net895 net3755 net412 VGND VGND VPWR VPWR _00852_ sky130_fd_sc_hd__mux2_1
XFILLER_107_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08049_ data_array.data1\[0\]\[55\] net1343 net1249 data_array.data1\[3\]\[55\] _05234_
+ VGND VGND VPWR VPWR _05235_ sky130_fd_sc_hd__a221o_1
XFILLER_123_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold960 tag_array.tag1\[2\]\[14\] VGND VGND VPWR VPWR net2611 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold971 tag_array.tag0\[4\]\[21\] VGND VGND VPWR VPWR net2622 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold982 data_array.data1\[4\]\[25\] VGND VGND VPWR VPWR net2633 sky130_fd_sc_hd__dlygate4sd3_1
X_11060_ net1764 net1020 net329 VGND VGND VPWR VPWR _02803_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_168_3581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold993 tag_array.tag1\[13\]\[21\] VGND VGND VPWR VPWR net2644 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_168_3592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10011_ net1041 net2170 net555 VGND VGND VPWR VPWR _01760_ sky130_fd_sc_hd__mux2_1
XFILLER_1_679 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_224_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_224_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_49_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_129_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2350 data_array.data0\[6\]\[10\] VGND VGND VPWR VPWR net4001 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2361 data_array.data0\[11\]\[39\] VGND VGND VPWR VPWR net4012 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2372 data_array.data1\[7\]\[52\] VGND VGND VPWR VPWR net4023 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2383 tag_array.tag1\[9\]\[3\] VGND VGND VPWR VPWR net4034 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2394 data_array.data0\[11\]\[37\] VGND VGND VPWR VPWR net4045 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1660 data_array.data1\[15\]\[49\] VGND VGND VPWR VPWR net3311 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1671 data_array.data1\[15\]\[59\] VGND VGND VPWR VPWR net3322 sky130_fd_sc_hd__dlygate4sd3_1
X_11962_ clknet_leaf_114_clk _00770_ VGND VGND VPWR VPWR data_array.data0\[4\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1682 data_array.data1\[6\]\[9\] VGND VGND VPWR VPWR net3333 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1693 data_array.data0\[12\]\[59\] VGND VGND VPWR VPWR net3344 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_151_86 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13701_ clknet_leaf_202_clk _02330_ VGND VGND VPWR VPWR data_array.data1\[15\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
X_10913_ net1090 net2803 net529 VGND VGND VPWR VPWR _02658_ sky130_fd_sc_hd__mux2_1
XFILLER_71_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11893_ clknet_leaf_34_clk _00701_ VGND VGND VPWR VPWR data_array.data0\[5\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13632_ clknet_leaf_230_clk _02261_ VGND VGND VPWR VPWR data_array.data0\[9\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
X_10844_ net1110 net3278 net517 VGND VGND VPWR VPWR _02589_ sky130_fd_sc_hd__mux2_1
XFILLER_71_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13563_ clknet_leaf_115_clk _02192_ VGND VGND VPWR VPWR data_array.data1\[0\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10775_ net874 net3920 net496 VGND VGND VPWR VPWR _02520_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12514_ clknet_leaf_179_clk _01208_ VGND VGND VPWR VPWR lru_array.lru_mem\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_9_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13494_ clknet_leaf_35_clk _02124_ VGND VGND VPWR VPWR tag_array.dirty1\[9\] sky130_fd_sc_hd__dfxtp_1
X_12445_ clknet_leaf_226_clk _01139_ VGND VGND VPWR VPWR data_array.data0\[14\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_176_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12376_ clknet_leaf_211_clk _00053_ VGND VGND VPWR VPWR data_array.rdata0\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_125_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14115_ clknet_leaf_238_clk _02744_ VGND VGND VPWR VPWR data_array.data0\[1\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_91_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11327_ net984 net4191 net800 VGND VGND VPWR VPWR _03070_ sky130_fd_sc_hd__mux2_1
X_14046_ clknet_leaf_24_clk _02675_ VGND VGND VPWR VPWR data_array.data1\[6\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_11258_ net998 net4569 net676 VGND VGND VPWR VPWR _03001_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_215_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_215_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10209_ net970 net3154 net355 VGND VGND VPWR VPWR _01956_ sky130_fd_sc_hd__mux2_1
XFILLER_79_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11189_ net1017 net4623 net652 VGND VGND VPWR VPWR _02932_ sky130_fd_sc_hd__mux2_1
XFILLER_67_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05750_ _03263_ _03264_ _03265_ _03266_ VGND VGND VPWR VPWR _03267_ sky130_fd_sc_hd__or4_1
XFILLER_82_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05681_ net9 fsm.tag_out0\[10\] VGND VGND VPWR VPWR _03198_ sky130_fd_sc_hd__and2b_1
XFILLER_39_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07420_ data_array.data0\[8\]\[62\] net1415 net1321 data_array.data0\[11\]\[62\]
+ _04662_ VGND VGND VPWR VPWR _04663_ sky130_fd_sc_hd__a221o_1
XFILLER_90_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_1069 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07351_ net1217 _04595_ _04599_ net1169 VGND VGND VPWR VPWR _04601_ sky130_fd_sc_hd__a22o_1
XFILLER_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06302_ tag_array.tag0\[8\]\[10\] net1405 net1311 tag_array.tag0\[11\]\[10\] _03646_
+ VGND VGND VPWR VPWR _03647_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_63_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07282_ data_array.data0\[5\]\[49\] net1580 net1484 data_array.data0\[6\]\[49\] VGND
+ VGND VPWR VPWR _04538_ sky130_fd_sc_hd__a22o_1
X_06233_ tag_array.tag0\[5\]\[4\] net1561 net1465 tag_array.tag0\[6\]\[4\] VGND VGND
+ VPWR VPWR _03584_ sky130_fd_sc_hd__a22o_1
X_09021_ net2572 net940 net424 VGND VGND VPWR VPWR _00776_ sky130_fd_sc_hd__mux2_1
XFILLER_129_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06164_ tag_array.valid0\[0\] net1407 net1313 tag_array.valid0\[3\] _03520_ VGND
+ VGND VPWR VPWR _03521_ sky130_fd_sc_hd__a221o_1
XFILLER_85_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold201 data_array.data1\[8\]\[9\] VGND VGND VPWR VPWR net1852 sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 tag_array.tag1\[8\]\[11\] VGND VGND VPWR VPWR net1863 sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 data_array.data0\[1\]\[62\] VGND VGND VPWR VPWR net1874 sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 data_array.data1\[1\]\[59\] VGND VGND VPWR VPWR net1885 sky130_fd_sc_hd__dlygate4sd3_1
X_06095_ data_array.rdata0\[10\] net1141 net1119 data_array.rdata1\[10\] VGND VGND
+ VPWR VPWR net264 sky130_fd_sc_hd__a22o_1
Xhold245 data_array.data0\[4\]\[36\] VGND VGND VPWR VPWR net1896 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold256 data_array.data1\[4\]\[44\] VGND VGND VPWR VPWR net1907 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold267 data_array.data0\[8\]\[29\] VGND VGND VPWR VPWR net1918 sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 data_array.data0\[0\]\[22\] VGND VGND VPWR VPWR net1929 sky130_fd_sc_hd__dlygate4sd3_1
X_09923_ net716 net3439 net603 VGND VGND VPWR VPWR _01673_ sky130_fd_sc_hd__mux2_1
Xfanout703 _05409_ VGND VGND VPWR VPWR net703 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold289 tag_array.tag1\[4\]\[2\] VGND VGND VPWR VPWR net1940 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout714 net717 VGND VGND VPWR VPWR net714 sky130_fd_sc_hd__clkbuf_2
Xfanout725 _05399_ VGND VGND VPWR VPWR net725 sky130_fd_sc_hd__buf_1
Xclkbuf_leaf_206_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_206_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_86_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout736 net737 VGND VGND VPWR VPWR net736 sky130_fd_sc_hd__clkbuf_2
Xfanout747 _05387_ VGND VGND VPWR VPWR net747 sky130_fd_sc_hd__buf_1
X_09854_ net1053 net3504 net382 VGND VGND VPWR VPWR _01604_ sky130_fd_sc_hd__mux2_1
XFILLER_59_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_24 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout758 net759 VGND VGND VPWR VPWR net758 sky130_fd_sc_hd__clkbuf_2
Xfanout769 _05377_ VGND VGND VPWR VPWR net769 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_146_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08805_ net2929 net1026 net444 VGND VGND VPWR VPWR _00563_ sky130_fd_sc_hd__mux2_1
XFILLER_100_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09785_ net1068 net2792 net392 VGND VGND VPWR VPWR _01536_ sky130_fd_sc_hd__mux2_1
X_06997_ data_array.data0\[4\]\[23\] net1366 net1272 data_array.data0\[7\]\[23\] _04278_
+ VGND VGND VPWR VPWR _04279_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_107_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08736_ net778 net3147 net457 VGND VGND VPWR VPWR _00495_ sky130_fd_sc_hd__mux2_1
XFILLER_73_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05948_ data_array.rdata0\[39\] net847 net1143 VGND VGND VPWR VPWR _03426_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_124_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08667_ net756 net4413 net500 VGND VGND VPWR VPWR _00426_ sky130_fd_sc_hd__mux2_1
X_05879_ data_array.rdata0\[16\] net848 net1144 VGND VGND VPWR VPWR _03380_ sky130_fd_sc_hd__o21a_1
XFILLER_42_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07618_ data_array.data1\[8\]\[16\] net1354 net1260 data_array.data1\[11\]\[16\]
+ _04842_ VGND VGND VPWR VPWR _04843_ sky130_fd_sc_hd__a221o_1
X_08598_ net730 net3387 net534 VGND VGND VPWR VPWR _00357_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_120_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07549_ net1178 _04775_ _04779_ net1226 VGND VGND VPWR VPWR _04781_ sky130_fd_sc_hd__a22o_1
X_10560_ net966 net3266 net461 VGND VGND VPWR VPWR _02305_ sky130_fd_sc_hd__mux2_1
XFILLER_14_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09219_ net704 net2588 net632 VGND VGND VPWR VPWR _00973_ sky130_fd_sc_hd__mux2_1
X_10491_ net982 net4222 net344 VGND VGND VPWR VPWR _02236_ sky130_fd_sc_hd__mux2_1
XFILLER_10_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_101_Left_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12230_ clknet_leaf_151_clk _00159_ VGND VGND VPWR VPWR fsm.tag_out1\[12\] sky130_fd_sc_hd__dfxtp_2
XFILLER_154_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_80_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12161_ clknet_leaf_181_clk _00969_ VGND VGND VPWR VPWR tag_array.tag0\[13\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_123_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11112_ net1071 net2940 net551 VGND VGND VPWR VPWR _02855_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12092_ clknet_leaf_77_clk _00900_ VGND VGND VPWR VPWR data_array.data1\[14\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_9_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold790 data_array.data0\[14\]\[46\] VGND VGND VPWR VPWR net2441 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11043_ net1911 net1089 net330 VGND VGND VPWR VPWR _02786_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_183_3876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2180 data_array.data1\[14\]\[52\] VGND VGND VPWR VPWR net3831 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_4_3_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_3_0_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_110_Left_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2191 data_array.data0\[15\]\[16\] VGND VGND VPWR VPWR net3842 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_64_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12994_ clknet_leaf_61_clk _01688_ VGND VGND VPWR VPWR data_array.data0\[3\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_91_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1490 tag_array.tag0\[8\]\[12\] VGND VGND VPWR VPWR net3141 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11945_ clknet_leaf_59_clk _00753_ VGND VGND VPWR VPWR data_array.data0\[4\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_55_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11876_ clknet_leaf_49_clk _00684_ VGND VGND VPWR VPWR data_array.data0\[5\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_177_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13615_ clknet_leaf_124_clk _02244_ VGND VGND VPWR VPWR data_array.data0\[9\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
X_10827_ net1790 net922 net509 VGND VGND VPWR VPWR _02572_ sky130_fd_sc_hd__mux2_1
XFILLER_158_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_1080 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13546_ clknet_leaf_36_clk _02175_ VGND VGND VPWR VPWR data_array.data1\[0\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
X_10758_ net942 net4471 net498 VGND VGND VPWR VPWR _02503_ sky130_fd_sc_hd__mux2_1
X_13477_ clknet_leaf_145_clk _02107_ VGND VGND VPWR VPWR tag_array.tag0\[15\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_10689_ net2465 net960 net481 VGND VGND VPWR VPWR _02434_ sky130_fd_sc_hd__mux2_1
X_12428_ clknet_leaf_22_clk _01122_ VGND VGND VPWR VPWR data_array.data0\[14\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_127_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput306 net306 VGND VGND VPWR VPWR mem_wdata[49] sky130_fd_sc_hd__buf_2
Xoutput317 net317 VGND VGND VPWR VPWR mem_wdata[59] sky130_fd_sc_hd__buf_2
XFILLER_99_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12359_ clknet_leaf_256_clk _00035_ VGND VGND VPWR VPWR data_array.rdata0\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_141_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14029_ clknet_leaf_201_clk _02658_ VGND VGND VPWR VPWR data_array.data1\[6\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_06920_ data_array.data0\[0\]\[16\] net1358 net1264 data_array.data0\[3\]\[16\] _04208_
+ VGND VGND VPWR VPWR _04209_ sky130_fd_sc_hd__a221o_1
XFILLER_67_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06851_ data_array.data0\[13\]\[10\] net1601 net1505 data_array.data0\[14\]\[10\]
+ VGND VGND VPWR VPWR _04146_ sky130_fd_sc_hd__a22o_1
XFILLER_83_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05802_ _03172_ _03183_ _03204_ net1654 VGND VGND VPWR VPWR _03319_ sky130_fd_sc_hd__or4_1
X_09570_ net1068 net2409 net400 VGND VGND VPWR VPWR _01322_ sky130_fd_sc_hd__mux2_1
X_06782_ data_array.data0\[8\]\[4\] net1391 net1297 data_array.data0\[11\]\[4\] _04082_
+ VGND VGND VPWR VPWR _04083_ sky130_fd_sc_hd__a221o_1
X_08521_ net1717 net599 VGND VGND VPWR VPWR _00301_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_141_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05733_ net6 fsm.tag_out1\[7\] VGND VGND VPWR VPWR _03250_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_141_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_65_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08452_ net1128 _05537_ VGND VGND VPWR VPWR _05538_ sky130_fd_sc_hd__and2_1
XFILLER_23_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05664_ _03178_ _03179_ _03180_ VGND VGND VPWR VPWR _03181_ sky130_fd_sc_hd__or3_1
XFILLER_51_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07403_ data_array.data0\[1\]\[60\] net1603 net1507 data_array.data0\[2\]\[60\] VGND
+ VGND VPWR VPWR _04648_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_82_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08383_ net1129 _05491_ VGND VGND VPWR VPWR _05492_ sky130_fd_sc_hd__and2_1
XFILLER_91_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_1014 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07334_ data_array.data0\[0\]\[54\] net1356 net1262 data_array.data0\[3\]\[54\] _04584_
+ VGND VGND VPWR VPWR _04585_ sky130_fd_sc_hd__a221o_1
XFILLER_177_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07265_ data_array.data0\[9\]\[48\] net1581 net1485 data_array.data0\[10\]\[48\]
+ VGND VGND VPWR VPWR _04522_ sky130_fd_sc_hd__a22o_1
XFILLER_176_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09004_ net2326 net1009 net418 VGND VGND VPWR VPWR _00759_ sky130_fd_sc_hd__mux2_1
X_06216_ tag_array.tag0\[0\]\[2\] net1368 net1274 tag_array.tag0\[3\]\[2\] _03568_
+ VGND VGND VPWR VPWR _03569_ sky130_fd_sc_hd__a221o_1
XFILLER_136_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07196_ net1616 _04453_ _04457_ net1190 VGND VGND VPWR VPWR _04460_ sky130_fd_sc_hd__a22o_1
X_06147_ data_array.rdata0\[62\] net1141 net1119 data_array.rdata1\[62\] VGND VGND
+ VPWR VPWR net321 sky130_fd_sc_hd__a22o_1
XFILLER_160_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_148_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_148_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06078_ fsm.tag_out0\[21\] net1122 _03502_ VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__a21o_1
Xfanout500 net501 VGND VGND VPWR VPWR net500 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_165_3540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1509 net1510 VGND VGND VPWR VPWR net1509 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout511 net512 VGND VGND VPWR VPWR net511 sky130_fd_sc_hd__clkbuf_8
X_09906_ net785 net4298 net602 VGND VGND VPWR VPWR _01656_ sky130_fd_sc_hd__mux2_1
Xfanout522 _05599_ VGND VGND VPWR VPWR net522 sky130_fd_sc_hd__clkbuf_4
Xfanout533 net534 VGND VGND VPWR VPWR net533 sky130_fd_sc_hd__buf_2
XFILLER_120_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout544 net547 VGND VGND VPWR VPWR net544 sky130_fd_sc_hd__buf_2
Xfanout555 net560 VGND VGND VPWR VPWR net555 sky130_fd_sc_hd__buf_4
Xfanout566 net572 VGND VGND VPWR VPWR net566 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_126_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09837_ net860 net2361 net393 VGND VGND VPWR VPWR _01588_ sky130_fd_sc_hd__mux2_1
Xfanout577 _05592_ VGND VGND VPWR VPWR net577 sky130_fd_sc_hd__clkbuf_4
XFILLER_58_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout588 net589 VGND VGND VPWR VPWR net588 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_161_3448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout599 net601 VGND VGND VPWR VPWR net599 sky130_fd_sc_hd__buf_4
XFILLER_100_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09768_ net1840 net715 net672 VGND VGND VPWR VPWR _01520_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_122_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08719_ net2207 net746 net474 VGND VGND VPWR VPWR _00478_ sky130_fd_sc_hd__mux2_1
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09699_ net793 net3079 net610 VGND VGND VPWR VPWR _01451_ sky130_fd_sc_hd__mux2_1
X_11730_ clknet_leaf_155_clk _00538_ VGND VGND VPWR VPWR tag_array.tag0\[9\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_155_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ clknet_leaf_31_clk _00469_ VGND VGND VPWR VPWR tag_array.tag1\[1\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_25_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13400_ clknet_leaf_131_clk _02030_ VGND VGND VPWR VPWR data_array.data1\[8\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_41_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10612_ net3930 net1015 net473 VGND VGND VPWR VPWR _02357_ sky130_fd_sc_hd__mux2_1
X_14380_ clknet_leaf_67_clk _03003_ VGND VGND VPWR VPWR data_array.data1\[10\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_179_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11592_ clknet_leaf_139_clk _00400_ VGND VGND VPWR VPWR tag_array.tag1\[4\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13331_ clknet_leaf_124_clk _01961_ VGND VGND VPWR VPWR data_array.data0\[10\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_823 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10543_ net1035 net2823 net461 VGND VGND VPWR VPWR _02288_ sky130_fd_sc_hd__mux2_1
XFILLER_167_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13262_ clknet_leaf_243_clk _01892_ VGND VGND VPWR VPWR data_array.data0\[11\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_108_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10474_ net1049 net3788 net349 VGND VGND VPWR VPWR _02219_ sky130_fd_sc_hd__mux2_1
XFILLER_183_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12213_ clknet_leaf_183_clk _00143_ VGND VGND VPWR VPWR fsm.tag_out0\[20\] sky130_fd_sc_hd__dfxtp_2
XFILLER_109_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13193_ clknet_leaf_68_clk _00087_ VGND VGND VPWR VPWR data_array.rdata1\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_29_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12144_ clknet_leaf_171_clk _00952_ VGND VGND VPWR VPWR tag_array.tag0\[13\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_111_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12075_ clknet_leaf_229_clk _00883_ VGND VGND VPWR VPWR data_array.data1\[14\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_11026_ net1886 net896 net336 VGND VGND VPWR VPWR _02770_ sky130_fd_sc_hd__mux2_1
XFILLER_65_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12977_ clknet_leaf_108_clk _01671_ VGND VGND VPWR VPWR tag_array.tag0\[4\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_92_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11928_ clknet_leaf_247_clk _00736_ VGND VGND VPWR VPWR data_array.data0\[4\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11859_ clknet_leaf_207_clk _00667_ VGND VGND VPWR VPWR data_array.data0\[7\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_18 _03477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_29 _05417_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13529_ clknet_leaf_254_clk _02158_ VGND VGND VPWR VPWR data_array.data1\[0\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_07050_ data_array.data0\[12\]\[28\] net1351 net1257 data_array.data0\[15\]\[28\]
+ _04326_ VGND VGND VPWR VPWR _04327_ sky130_fd_sc_hd__a221o_1
XFILLER_174_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06001_ net150 net1154 _03460_ _03461_ VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__a22o_1
XFILLER_127_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput169 net169 VGND VGND VPWR VPWR cpu_rdata[13] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_58_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2905 tag_array.dirty1\[5\] VGND VGND VPWR VPWR net4556 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_99_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07952_ data_array.data1\[12\]\[46\] net1333 net1239 data_array.data1\[15\]\[46\]
+ _05146_ VGND VGND VPWR VPWR _05147_ sky130_fd_sc_hd__a221o_1
XFILLER_102_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2916 tag_array.tag1\[6\]\[9\] VGND VGND VPWR VPWR net4567 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2927 data_array.data1\[7\]\[53\] VGND VGND VPWR VPWR net4578 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2938 data_array.data1\[11\]\[39\] VGND VGND VPWR VPWR net4589 sky130_fd_sc_hd__dlygate4sd3_1
X_06903_ data_array.data0\[8\]\[15\] net1394 net1300 data_array.data0\[11\]\[15\]
+ _04192_ VGND VGND VPWR VPWR _04193_ sky130_fd_sc_hd__a221o_1
Xhold2949 data_array.data1\[5\]\[61\] VGND VGND VPWR VPWR net4600 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_68_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_143_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07883_ data_array.data1\[5\]\[40\] net1605 net1509 data_array.data1\[6\]\[40\] VGND
+ VGND VPWR VPWR _05084_ sky130_fd_sc_hd__a22o_1
XFILLER_110_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09622_ net860 net2261 net401 VGND VGND VPWR VPWR _01374_ sky130_fd_sc_hd__mux2_1
XFILLER_68_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06834_ net1168 _04125_ _04129_ net1216 VGND VGND VPWR VPWR _04131_ sky130_fd_sc_hd__a22o_1
XFILLER_95_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09553_ net716 net2677 net619 VGND VGND VPWR VPWR _01306_ sky130_fd_sc_hd__mux2_1
X_06765_ data_array.data0\[1\]\[2\] net1528 net1432 data_array.data0\[2\]\[2\] VGND
+ VGND VPWR VPWR _04068_ sky130_fd_sc_hd__a22o_1
XFILLER_71_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08504_ net824 net813 _05361_ net855 VGND VGND VPWR VPWR _05573_ sky130_fd_sc_hd__or4_1
X_05716_ _03174_ _03175_ _03195_ _03208_ VGND VGND VPWR VPWR _03233_ sky130_fd_sc_hd__or4_1
XFILLER_24_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09484_ net794 net2776 net625 VGND VGND VPWR VPWR _01237_ sky130_fd_sc_hd__mux2_1
X_06696_ tag_array.tag1\[4\]\[21\] net1403 net1309 tag_array.tag1\[7\]\[21\] _04004_
+ VGND VGND VPWR VPWR _04005_ sky130_fd_sc_hd__a221o_1
XFILLER_51_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08435_ net2151 net896 net686 VGND VGND VPWR VPWR _00274_ sky130_fd_sc_hd__mux2_1
XFILLER_52_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05647_ net32 fsm.tag_out0\[2\] VGND VGND VPWR VPWR _03164_ sky130_fd_sc_hd__nand2_1
XFILLER_178_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08366_ net2081 net989 net691 VGND VGND VPWR VPWR _00251_ sky130_fd_sc_hd__mux2_1
X_07317_ net1195 _04563_ _04567_ net1621 VGND VGND VPWR VPWR _04570_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_119_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08297_ net2711 net1080 net693 VGND VGND VPWR VPWR _00228_ sky130_fd_sc_hd__mux2_1
XFILLER_178_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07248_ data_array.data0\[12\]\[46\] net1341 net1247 data_array.data0\[15\]\[46\]
+ _04506_ VGND VGND VPWR VPWR _04507_ sky130_fd_sc_hd__a221o_1
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07179_ data_array.data0\[5\]\[40\] net1602 net1506 data_array.data0\[6\]\[40\] VGND
+ VGND VPWR VPWR _04444_ sky130_fd_sc_hd__a22o_1
XFILLER_180_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10190_ net1046 net4232 net356 VGND VGND VPWR VPWR _01937_ sky130_fd_sc_hd__mux2_1
XFILLER_160_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1306 _03515_ VGND VGND VPWR VPWR net1306 sky130_fd_sc_hd__buf_4
XFILLER_105_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1317 net1319 VGND VGND VPWR VPWR net1317 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_180_3813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout330 net331 VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__buf_4
Xfanout1328 _03515_ VGND VGND VPWR VPWR net1328 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_180_3824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1339 net1376 VGND VGND VPWR VPWR net1339 sky130_fd_sc_hd__buf_2
Xfanout341 net342 VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__buf_4
Xfanout352 _03130_ VGND VGND VPWR VPWR net352 sky130_fd_sc_hd__clkbuf_2
XFILLER_120_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout363 net369 VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__clkbuf_8
XFILLER_115_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout374 _03127_ VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__clkbuf_4
Xfanout385 _03126_ VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__buf_4
XFILLER_87_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12900_ clknet_leaf_71_clk _01594_ VGND VGND VPWR VPWR data_array.data0\[13\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout396 net397 VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__buf_4
XFILLER_47_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13880_ clknet_leaf_75_clk _02509_ VGND VGND VPWR VPWR data_array.data1\[3\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_143_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12831_ clknet_leaf_188_clk _01525_ VGND VGND VPWR VPWR tag_array.tag1\[0\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12762_ clknet_leaf_143_clk _01456_ VGND VGND VPWR VPWR tag_array.tag0\[6\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_178_3775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_3786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14501_ clknet_leaf_175_clk _03122_ VGND VGND VPWR VPWR lru_array.lru_mem\[5\] sky130_fd_sc_hd__dfxtp_1
X_11713_ clknet_leaf_178_clk _00521_ VGND VGND VPWR VPWR tag_array.tag0\[9\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12693_ clknet_leaf_161_clk _01387_ VGND VGND VPWR VPWR tag_array.tag0\[8\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14432_ clknet_leaf_212_clk _03055_ VGND VGND VPWR VPWR data_array.data1\[7\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_11644_ clknet_leaf_102_clk _00452_ VGND VGND VPWR VPWR tag_array.tag1\[2\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_155_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14363_ clknet_leaf_199_clk _02986_ VGND VGND VPWR VPWR data_array.data1\[10\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_11575_ clknet_leaf_140_clk _00383_ VGND VGND VPWR VPWR tag_array.tag1\[5\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput16 cpu_addr[23] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput27 cpu_addr[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_4
Xinput38 cpu_wdata[13] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_1
X_13314_ clknet_leaf_176_clk _01944_ VGND VGND VPWR VPWR data_array.data0\[10\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_10526_ net1101 net3570 net454 VGND VGND VPWR VPWR _02271_ sky130_fd_sc_hd__mux2_1
Xinput49 cpu_wdata[23] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_1
XFILLER_182_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14294_ clknet_leaf_42_clk _02923_ VGND VGND VPWR VPWR data_array.data1\[11\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_155_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13245_ clknet_leaf_16_clk _01875_ VGND VGND VPWR VPWR data_array.data0\[11\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_170_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10457_ net353 net4049 net456 VGND VGND VPWR VPWR _02203_ sky130_fd_sc_hd__mux2_1
XFILLER_124_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13176_ clknet_leaf_201_clk _00068_ VGND VGND VPWR VPWR data_array.rdata1\[13\] sky130_fd_sc_hd__dfxtp_1
X_10388_ net1829 net1100 net661 VGND VGND VPWR VPWR _02134_ sky130_fd_sc_hd__mux2_1
XFILLER_151_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12127_ clknet_leaf_158_clk _00935_ VGND VGND VPWR VPWR tag_array.tag0\[12\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_12058_ clknet_leaf_68_clk _00866_ VGND VGND VPWR VPWR data_array.data1\[14\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11009_ net2220 net964 net343 VGND VGND VPWR VPWR _02753_ sky130_fd_sc_hd__mux2_1
XFILLER_77_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06550_ tag_array.tag1\[9\]\[8\] net1608 net1512 tag_array.tag1\[10\]\[8\] VGND VGND
+ VPWR VPWR _03872_ sky130_fd_sc_hd__a22o_1
XFILLER_80_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06481_ net1199 _03803_ _03807_ net1625 VGND VGND VPWR VPWR _03810_ sky130_fd_sc_hd__a22o_1
XFILLER_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08220_ net759 net3242 net805 VGND VGND VPWR VPWR _00204_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08151_ tag_array.dirty1\[5\] net1540 net1444 tag_array.dirty1\[6\] VGND VGND VPWR
+ VPWR _05328_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_99_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07102_ data_array.data0\[1\]\[33\] net1585 net1489 data_array.data0\[2\]\[33\] VGND
+ VGND VPWR VPWR _04374_ sky130_fd_sc_hd__a22o_1
Xclkload210 clknet_leaf_117_clk VGND VGND VPWR VPWR clkload210/Y sky130_fd_sc_hd__inv_8
X_08082_ data_array.data1\[4\]\[58\] net1359 net1265 data_array.data1\[7\]\[58\] _05264_
+ VGND VGND VPWR VPWR _05265_ sky130_fd_sc_hd__a221o_1
Xclkload221 clknet_leaf_156_clk VGND VGND VPWR VPWR clkload221/Y sky130_fd_sc_hd__clkinv_4
Xclkload232 clknet_leaf_130_clk VGND VGND VPWR VPWR clkload232/Y sky130_fd_sc_hd__clkinv_4
Xclkload243 clknet_leaf_140_clk VGND VGND VPWR VPWR clkload243/Y sky130_fd_sc_hd__clkinv_4
XFILLER_161_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07033_ _04310_ _04311_ VGND VGND VPWR VPWR _00018_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_77_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08984_ net1877 net1088 net420 VGND VGND VPWR VPWR _00739_ sky130_fd_sc_hd__mux2_1
XFILLER_87_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2702 data_array.data1\[3\]\[29\] VGND VGND VPWR VPWR net4353 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2713 data_array.data1\[5\]\[5\] VGND VGND VPWR VPWR net4364 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2724 data_array.data0\[14\]\[27\] VGND VGND VPWR VPWR net4375 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_110_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2735 tag_array.tag1\[11\]\[14\] VGND VGND VPWR VPWR net4386 sky130_fd_sc_hd__dlygate4sd3_1
X_07935_ _05130_ _05131_ VGND VGND VPWR VPWR _00102_ sky130_fd_sc_hd__or2_1
Xhold2746 data_array.data1\[14\]\[54\] VGND VGND VPWR VPWR net4397 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2757 tag_array.tag0\[11\]\[7\] VGND VGND VPWR VPWR net4408 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2768 tag_array.tag1\[10\]\[13\] VGND VGND VPWR VPWR net4419 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2779 tag_array.tag1\[15\]\[19\] VGND VGND VPWR VPWR net4430 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07866_ data_array.data1\[4\]\[38\] net1397 net1303 data_array.data1\[7\]\[38\] _05068_
+ VGND VGND VPWR VPWR _05069_ sky130_fd_sc_hd__a221o_1
XFILLER_29_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09605_ net928 net3685 net395 VGND VGND VPWR VPWR _01357_ sky130_fd_sc_hd__mux2_1
XFILLER_83_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06817_ data_array.data0\[0\]\[7\] net1411 net1317 data_array.data0\[3\]\[7\] _04114_
+ VGND VGND VPWR VPWR _04115_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_27_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07797_ data_array.data1\[9\]\[32\] net1520 net1424 data_array.data1\[10\]\[32\]
+ VGND VGND VPWR VPWR _05006_ sky130_fd_sc_hd__a22o_1
XFILLER_84_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09536_ net784 net4118 net618 VGND VGND VPWR VPWR _01289_ sky130_fd_sc_hd__mux2_1
X_06748_ data_array.data0\[13\]\[1\] net1523 net1427 data_array.data0\[14\]\[1\] VGND
+ VGND VPWR VPWR _04052_ sky130_fd_sc_hd__a22o_1
XFILLER_58_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09467_ net760 net2314 net659 VGND VGND VPWR VPWR _01220_ sky130_fd_sc_hd__mux2_1
X_06679_ net1634 _03983_ _03987_ net1208 VGND VGND VPWR VPWR _03990_ sky130_fd_sc_hd__a22o_1
XFILLER_40_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08418_ net141 net76 net1642 VGND VGND VPWR VPWR _05515_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_156_3358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09398_ net1075 net2815 net586 VGND VGND VPWR VPWR _01151_ sky130_fd_sc_hd__mux2_1
XFILLER_145_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_3683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08349_ net116 net51 net1638 VGND VGND VPWR VPWR _05469_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_117_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_173_3694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_129_Right_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11360_ net820 net2414 _05605_ VGND VGND VPWR VPWR _03103_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_134_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10311_ net2108 net919 net640 VGND VGND VPWR VPWR _02058_ sky130_fd_sc_hd__mux2_1
XFILLER_4_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11291_ net864 net3271 net677 VGND VGND VPWR VPWR _03034_ sky130_fd_sc_hd__mux2_1
XFILLER_3_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13030_ clknet_leaf_20_clk _01724_ VGND VGND VPWR VPWR data_array.data0\[3\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
X_10242_ net776 net3104 net595 VGND VGND VPWR VPWR _01989_ sky130_fd_sc_hd__mux2_1
XFILLER_3_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1103 _05424_ VGND VGND VPWR VPWR net1103 sky130_fd_sc_hd__buf_1
X_10173_ net807 _05547_ VGND VGND VPWR VPWR _03129_ sky130_fd_sc_hd__nand2_1
XFILLER_105_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1114 net1115 VGND VGND VPWR VPWR net1114 sky130_fd_sc_hd__clkbuf_4
Xfanout1125 net1130 VGND VGND VPWR VPWR net1125 sky130_fd_sc_hd__clkbuf_4
Xfanout1136 net1137 VGND VGND VPWR VPWR net1136 sky130_fd_sc_hd__clkbuf_4
Xfanout1147 net1148 VGND VGND VPWR VPWR net1147 sky130_fd_sc_hd__buf_4
XFILLER_154_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1158 net1160 VGND VGND VPWR VPWR net1158 sky130_fd_sc_hd__buf_2
Xfanout1169 net1175 VGND VGND VPWR VPWR net1169 sky130_fd_sc_hd__buf_4
XFILLER_87_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13932_ clknet_leaf_117_clk _02561_ VGND VGND VPWR VPWR data_array.data1\[4\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13863_ clknet_leaf_41_clk _02492_ VGND VGND VPWR VPWR data_array.data1\[3\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12814_ clknet_leaf_132_clk _01508_ VGND VGND VPWR VPWR tag_array.tag1\[0\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13794_ clknet_leaf_255_clk _02423_ VGND VGND VPWR VPWR data_array.data1\[2\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_5_21__f_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_5_21__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_12745_ clknet_leaf_146_clk _01439_ VGND VGND VPWR VPWR tag_array.tag0\[5\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12676_ clknet_leaf_207_clk _01370_ VGND VGND VPWR VPWR data_array.data0\[15\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_13_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14415_ clknet_leaf_172_clk _03038_ VGND VGND VPWR VPWR lru_array.lru_mem\[14\] sky130_fd_sc_hd__dfxtp_1
X_11627_ clknet_leaf_187_clk _00435_ VGND VGND VPWR VPWR tag_array.tag1\[3\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_14346_ clknet_leaf_185_clk _00183_ _00191_ VGND VGND VPWR VPWR fsm.state\[2\] sky130_fd_sc_hd__dfrtp_4
X_11558_ clknet_leaf_189_clk _00366_ VGND VGND VPWR VPWR tag_array.tag1\[6\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold608 data_array.data1\[8\]\[16\] VGND VGND VPWR VPWR net2259 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10509_ net910 net3591 net351 VGND VGND VPWR VPWR _02254_ sky130_fd_sc_hd__mux2_1
X_14277_ clknet_leaf_203_clk _02906_ VGND VGND VPWR VPWR data_array.data1\[12\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold619 tag_array.tag1\[0\]\[11\] VGND VGND VPWR VPWR net2270 sky130_fd_sc_hd__dlygate4sd3_1
X_11489_ clknet_leaf_155_clk _00298_ VGND VGND VPWR VPWR tag_array.valid0\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_94_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13228_ clknet_leaf_5_clk _01858_ VGND VGND VPWR VPWR data_array.data0\[11\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_171_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13159_ clknet_leaf_101_clk _01853_ VGND VGND VPWR VPWR tag_array.tag1\[8\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2009 tag_array.tag0\[3\]\[19\] VGND VGND VPWR VPWR net3660 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_98_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05981_ data_array.rdata0\[50\] net846 net1143 VGND VGND VPWR VPWR _03448_ sky130_fd_sc_hd__o21a_1
Xhold1308 data_array.data0\[7\]\[24\] VGND VGND VPWR VPWR net2959 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1319 data_array.data0\[3\]\[40\] VGND VGND VPWR VPWR net2970 sky130_fd_sc_hd__dlygate4sd3_1
X_07720_ data_array.data1\[9\]\[25\] net1520 net1424 data_array.data1\[10\]\[25\]
+ VGND VGND VPWR VPWR _04936_ sky130_fd_sc_hd__a22o_1
XFILLER_77_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07651_ data_array.data1\[12\]\[19\] net1394 net1300 data_array.data1\[15\]\[19\]
+ _04872_ VGND VGND VPWR VPWR _04873_ sky130_fd_sc_hd__a221o_1
XFILLER_81_802 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06602_ net1207 _03913_ _03917_ net1633 VGND VGND VPWR VPWR _03920_ sky130_fd_sc_hd__a22o_1
XFILLER_92_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07582_ net1231 _04805_ _04809_ net1179 VGND VGND VPWR VPWR _04811_ sky130_fd_sc_hd__a22o_1
X_09321_ net695 net3611 net546 VGND VGND VPWR VPWR _01075_ sky130_fd_sc_hd__mux2_1
X_06533_ tag_array.tag1\[8\]\[6\] net1362 net1268 tag_array.tag1\[11\]\[6\] _03856_
+ VGND VGND VPWR VPWR _03857_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_138_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09252_ net772 net3451 net576 VGND VGND VPWR VPWR _01006_ sky130_fd_sc_hd__mux2_1
XFILLER_22_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06464_ tag_array.tag1\[1\]\[0\] net1576 net1480 tag_array.tag1\[2\]\[0\] VGND VGND
+ VPWR VPWR _03794_ sky130_fd_sc_hd__a22o_1
XFILLER_22_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08203_ net1649 net1158 net2 VGND VGND VPWR VPWR _05370_ sky130_fd_sc_hd__and3_1
X_09183_ net748 net2877 net627 VGND VGND VPWR VPWR _00937_ sky130_fd_sc_hd__mux2_1
XFILLER_21_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06395_ _03730_ _03731_ VGND VGND VPWR VPWR _00140_ sky130_fd_sc_hd__or2_1
XFILLER_175_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08134_ data_array.data1\[13\]\[63\] net1553 net1457 data_array.data1\[14\]\[63\]
+ VGND VGND VPWR VPWR _05312_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_151_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_612 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08065_ net1192 _05243_ _05247_ net1618 VGND VGND VPWR VPWR _05250_ sky130_fd_sc_hd__a22o_1
XFILLER_88_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_1027 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07016_ data_array.data0\[9\]\[25\] net1522 net1426 data_array.data0\[10\]\[25\]
+ VGND VGND VPWR VPWR _04296_ sky130_fd_sc_hd__a22o_1
XFILLER_150_829 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_712 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2510 data_array.data1\[10\]\[4\] VGND VGND VPWR VPWR net4161 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2521 data_array.data1\[3\]\[54\] VGND VGND VPWR VPWR net4172 sky130_fd_sc_hd__dlygate4sd3_1
X_08967_ net896 net3193 net426 VGND VGND VPWR VPWR _00723_ sky130_fd_sc_hd__mux2_1
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2532 tag_array.tag0\[4\]\[24\] VGND VGND VPWR VPWR net4183 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2543 tag_array.tag0\[4\]\[11\] VGND VGND VPWR VPWR net4194 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2554 data_array.data0\[6\]\[30\] VGND VGND VPWR VPWR net4205 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2565 data_array.data0\[6\]\[60\] VGND VGND VPWR VPWR net4216 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1820 data_array.data0\[9\]\[9\] VGND VGND VPWR VPWR net3471 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_25_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07918_ data_array.data1\[13\]\[43\] net1568 net1472 data_array.data1\[14\]\[43\]
+ VGND VGND VPWR VPWR _05116_ sky130_fd_sc_hd__a22o_1
Xhold1831 data_array.data0\[3\]\[59\] VGND VGND VPWR VPWR net3482 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2576 tag_array.tag0\[0\]\[13\] VGND VGND VPWR VPWR net4227 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1842 data_array.data0\[14\]\[16\] VGND VGND VPWR VPWR net3493 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08898_ net912 net3776 net438 VGND VGND VPWR VPWR _00655_ sky130_fd_sc_hd__mux2_1
Xhold2587 data_array.data0\[5\]\[44\] VGND VGND VPWR VPWR net4238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2598 data_array.data0\[15\]\[60\] VGND VGND VPWR VPWR net4249 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1853 data_array.data0\[13\]\[14\] VGND VGND VPWR VPWR net3504 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1864 tag_array.tag0\[6\]\[23\] VGND VGND VPWR VPWR net3515 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1875 tag_array.tag1\[11\]\[17\] VGND VGND VPWR VPWR net3526 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1886 data_array.data0\[9\]\[44\] VGND VGND VPWR VPWR net3537 sky130_fd_sc_hd__dlygate4sd3_1
X_07849_ data_array.data1\[8\]\[37\] net1353 net1259 data_array.data1\[11\]\[37\]
+ _05052_ VGND VGND VPWR VPWR _05053_ sky130_fd_sc_hd__a221o_1
XFILLER_72_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1897 tag_array.tag0\[6\]\[13\] VGND VGND VPWR VPWR net3548 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_158_3409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10860_ net1044 net3722 net516 VGND VGND VPWR VPWR _02605_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_175_3723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09519_ net752 net2709 net622 VGND VGND VPWR VPWR _01272_ sky130_fd_sc_hd__mux2_1
X_10791_ net1995 net1066 net507 VGND VGND VPWR VPWR _02536_ sky130_fd_sc_hd__mux2_1
XFILLER_40_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12530_ clknet_leaf_166_clk _01224_ VGND VGND VPWR VPWR tag_array.tag1\[11\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12461_ clknet_leaf_199_clk _01155_ VGND VGND VPWR VPWR data_array.data1\[9\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14200_ clknet_leaf_56_clk _02829_ VGND VGND VPWR VPWR data_array.data0\[2\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
X_11412_ clknet_leaf_262_clk _00222_ VGND VGND VPWR VPWR data_array.data0\[0\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_12392_ clknet_leaf_111_clk _01086_ VGND VGND VPWR VPWR data_array.data0\[14\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_153_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14131_ clknet_leaf_49_clk _02760_ VGND VGND VPWR VPWR data_array.data0\[1\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
X_11343_ net922 net3273 net802 VGND VGND VPWR VPWR _03086_ sky130_fd_sc_hd__mux2_1
XFILLER_181_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14062_ clknet_leaf_74_clk _02691_ VGND VGND VPWR VPWR data_array.data1\[6\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
X_11274_ net935 net4102 net682 VGND VGND VPWR VPWR _03017_ sky130_fd_sc_hd__mux2_1
XFILLER_3_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13013_ clknet_leaf_29_clk _01707_ VGND VGND VPWR VPWR data_array.data0\[3\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_10225_ net905 net3809 net354 VGND VGND VPWR VPWR _01972_ sky130_fd_sc_hd__mux2_1
XFILLER_133_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10156_ net920 net4115 net366 VGND VGND VPWR VPWR _01904_ sky130_fd_sc_hd__mux2_1
XFILLER_181_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10087_ net2359 net774 net638 VGND VGND VPWR VPWR _01836_ sky130_fd_sc_hd__mux2_1
X_13915_ clknet_leaf_66_clk _02544_ VGND VGND VPWR VPWR data_array.data1\[4\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13846_ clknet_leaf_46_clk _02475_ VGND VGND VPWR VPWR data_array.data1\[3\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13777_ clknet_leaf_58_clk _02406_ VGND VGND VPWR VPWR data_array.data1\[2\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_10989_ net2048 net1047 net338 VGND VGND VPWR VPWR _02733_ sky130_fd_sc_hd__mux2_1
XFILLER_128_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12728_ clknet_leaf_156_clk _01422_ VGND VGND VPWR VPWR tag_array.tag0\[7\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_12659_ clknet_leaf_260_clk _01353_ VGND VGND VPWR VPWR data_array.data0\[15\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_96_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_962 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06180_ tag_array.valid1\[9\] net1559 net1463 tag_array.valid1\[10\] VGND VGND VPWR
+ VPWR _03536_ sky130_fd_sc_hd__a22o_1
XFILLER_8_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14329_ clknet_leaf_56_clk _02958_ VGND VGND VPWR VPWR data_array.data1\[11\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold405 data_array.data0\[0\]\[4\] VGND VGND VPWR VPWR net2056 sky130_fd_sc_hd__dlygate4sd3_1
Xhold416 data_array.data0\[13\]\[19\] VGND VGND VPWR VPWR net2067 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold427 data_array.data0\[4\]\[37\] VGND VGND VPWR VPWR net2078 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold438 data_array.data0\[0\]\[24\] VGND VGND VPWR VPWR net2089 sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 data_array.data1\[0\]\[38\] VGND VGND VPWR VPWR net2100 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09870_ net989 net3320 net383 VGND VGND VPWR VPWR _01620_ sky130_fd_sc_hd__mux2_1
Xfanout907 _05522_ VGND VGND VPWR VPWR net907 sky130_fd_sc_hd__buf_1
Xfanout918 _05516_ VGND VGND VPWR VPWR net918 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_70_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout929 _05510_ VGND VGND VPWR VPWR net929 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_135_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08821_ net1899 net962 net444 VGND VGND VPWR VPWR _00579_ sky130_fd_sc_hd__mux2_1
Xhold1105 data_array.data1\[5\]\[50\] VGND VGND VPWR VPWR net2756 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1116 tag_array.tag1\[0\]\[14\] VGND VGND VPWR VPWR net2767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1127 tag_array.tag0\[12\]\[12\] VGND VGND VPWR VPWR net2778 sky130_fd_sc_hd__dlygate4sd3_1
X_08752_ net714 net4430 net460 VGND VGND VPWR VPWR _00511_ sky130_fd_sc_hd__mux2_1
X_05964_ data_array.rdata1\[44\] net834 net843 VGND VGND VPWR VPWR _03437_ sky130_fd_sc_hd__a21o_1
Xhold1138 data_array.data1\[4\]\[48\] VGND VGND VPWR VPWR net2789 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1149 data_array.data1\[14\]\[36\] VGND VGND VPWR VPWR net2800 sky130_fd_sc_hd__dlygate4sd3_1
X_07703_ net1219 _04915_ _04919_ net1171 VGND VGND VPWR VPWR _04921_ sky130_fd_sc_hd__a22o_1
XFILLER_38_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_876 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08683_ net2748 net791 net483 VGND VGND VPWR VPWR _00442_ sky130_fd_sc_hd__mux2_1
X_05895_ data_array.rdata1\[21\] net830 net839 VGND VGND VPWR VPWR _03391_ sky130_fd_sc_hd__a21o_1
X_07634_ data_array.data1\[5\]\[17\] net1526 net1430 data_array.data1\[6\]\[17\] VGND
+ VGND VPWR VPWR _04858_ sky130_fd_sc_hd__a22o_1
XFILLER_26_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_105_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07565_ data_array.data1\[0\]\[11\] net1384 net1290 data_array.data1\[3\]\[11\] _04794_
+ VGND VGND VPWR VPWR _04795_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_105_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_698 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09304_ net765 net2949 net551 VGND VGND VPWR VPWR _01058_ sky130_fd_sc_hd__mux2_1
XFILLER_55_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06516_ _03840_ _03841_ VGND VGND VPWR VPWR _00175_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_153_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07496_ data_array.data1\[9\]\[5\] net1551 net1455 data_array.data1\[10\]\[5\] VGND
+ VGND VPWR VPWR _04732_ sky130_fd_sc_hd__a22o_1
XFILLER_22_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09235_ net738 net3136 net646 VGND VGND VPWR VPWR _00989_ sky130_fd_sc_hd__mux2_1
XFILLER_142_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06447_ tag_array.tag0\[4\]\[23\] net1412 net1318 tag_array.tag0\[7\]\[23\] _03778_
+ VGND VGND VPWR VPWR _03779_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_170_3620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09166_ net879 net2291 net570 VGND VGND VPWR VPWR _00920_ sky130_fd_sc_hd__mux2_1
XFILLER_119_12 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06378_ tag_array.tag0\[9\]\[17\] net1602 net1506 tag_array.tag0\[10\]\[17\] VGND
+ VGND VPWR VPWR _03716_ sky130_fd_sc_hd__a22o_1
XFILLER_107_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08117_ data_array.data1\[8\]\[61\] net1354 net1260 data_array.data1\[11\]\[61\]
+ _05296_ VGND VGND VPWR VPWR _05297_ sky130_fd_sc_hd__a221o_1
XFILLER_163_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09097_ net896 net2738 net410 VGND VGND VPWR VPWR _00851_ sky130_fd_sc_hd__mux2_1
XFILLER_79_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08048_ data_array.data1\[1\]\[55\] net1534 net1438 data_array.data1\[2\]\[55\] VGND
+ VGND VPWR VPWR _05234_ sky130_fd_sc_hd__a22o_1
XFILLER_102_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold950 data_array.data0\[12\]\[36\] VGND VGND VPWR VPWR net2601 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold961 data_array.data0\[3\]\[62\] VGND VGND VPWR VPWR net2612 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_134_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold972 data_array.data0\[0\]\[44\] VGND VGND VPWR VPWR net2623 sky130_fd_sc_hd__dlygate4sd3_1
Xhold983 data_array.data1\[5\]\[2\] VGND VGND VPWR VPWR net2634 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_168_3582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold994 data_array.data1\[4\]\[55\] VGND VGND VPWR VPWR net2645 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_168_3593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10010_ net1045 net3834 net558 VGND VGND VPWR VPWR _01759_ sky130_fd_sc_hd__mux2_1
X_09999_ net1091 net3324 net558 VGND VGND VPWR VPWR _01748_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2340 tag_array.tag0\[10\]\[7\] VGND VGND VPWR VPWR net3991 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2351 data_array.data1\[11\]\[9\] VGND VGND VPWR VPWR net4002 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2362 data_array.data1\[13\]\[59\] VGND VGND VPWR VPWR net4013 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2373 data_array.data1\[14\]\[3\] VGND VGND VPWR VPWR net4024 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2384 tag_array.tag1\[11\]\[20\] VGND VGND VPWR VPWR net4035 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1650 data_array.data0\[11\]\[10\] VGND VGND VPWR VPWR net3301 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_971 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2395 data_array.data1\[7\]\[59\] VGND VGND VPWR VPWR net4046 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11961_ clknet_leaf_242_clk _00769_ VGND VGND VPWR VPWR data_array.data0\[4\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_57_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1661 data_array.data1\[11\]\[24\] VGND VGND VPWR VPWR net3312 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1672 data_array.data0\[5\]\[43\] VGND VGND VPWR VPWR net3323 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1683 data_array.data1\[2\]\[29\] VGND VGND VPWR VPWR net3334 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1694 data_array.data0\[5\]\[28\] VGND VGND VPWR VPWR net3345 sky130_fd_sc_hd__dlygate4sd3_1
X_13700_ clknet_leaf_119_clk _02329_ VGND VGND VPWR VPWR data_array.data1\[15\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_174_Left_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10912_ net1094 net4069 net532 VGND VGND VPWR VPWR _02657_ sky130_fd_sc_hd__mux2_1
XFILLER_72_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11892_ clknet_leaf_71_clk _00700_ VGND VGND VPWR VPWR data_array.data0\[5\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_13631_ clknet_leaf_12_clk _02260_ VGND VGND VPWR VPWR data_array.data0\[9\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
X_10843_ net1876 net858 net505 VGND VGND VPWR VPWR _02588_ sky130_fd_sc_hd__mux2_1
XFILLER_32_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13562_ clknet_leaf_41_clk _02191_ VGND VGND VPWR VPWR data_array.data1\[0\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
X_10774_ net878 net3795 net494 VGND VGND VPWR VPWR _02519_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_181_Right_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12513_ clknet_leaf_176_clk _01207_ VGND VGND VPWR VPWR lru_array.lru_mem\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_157_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13493_ clknet_leaf_182_clk _02123_ VGND VGND VPWR VPWR tag_array.tag0\[15\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_160_clk clknet_5_25__leaf_clk VGND VGND VPWR VPWR clknet_leaf_160_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_12_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12444_ clknet_leaf_110_clk _01138_ VGND VGND VPWR VPWR data_array.data0\[14\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_154_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_612 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_183_Left_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12375_ clknet_leaf_252_clk _00052_ VGND VGND VPWR VPWR data_array.rdata0\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_125_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14114_ clknet_leaf_246_clk _02743_ VGND VGND VPWR VPWR data_array.data0\[1\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_91_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11326_ net990 net3849 net801 VGND VGND VPWR VPWR _03069_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14045_ clknet_leaf_229_clk _02674_ VGND VGND VPWR VPWR data_array.data1\[6\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_180_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11257_ net1001 net2889 net674 VGND VGND VPWR VPWR _03000_ sky130_fd_sc_hd__mux2_1
XFILLER_79_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10208_ net972 net4330 net354 VGND VGND VPWR VPWR _01955_ sky130_fd_sc_hd__mux2_1
XFILLER_95_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11188_ net1021 net4594 net650 VGND VGND VPWR VPWR _02931_ sky130_fd_sc_hd__mux2_1
X_10139_ net989 net4508 net367 VGND VGND VPWR VPWR _01887_ sky130_fd_sc_hd__mux2_1
XFILLER_94_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05680_ _03193_ _03194_ _03195_ _03196_ VGND VGND VPWR VPWR _03197_ sky130_fd_sc_hd__or4_4
XFILLER_35_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13829_ clknet_leaf_211_clk _02458_ VGND VGND VPWR VPWR data_array.data1\[2\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_67_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07350_ net1192 _04593_ _04597_ net1618 VGND VGND VPWR VPWR _04600_ sky130_fd_sc_hd__a22o_1
X_06301_ tag_array.tag0\[9\]\[10\] net1602 net1506 tag_array.tag0\[10\]\[10\] VGND
+ VGND VPWR VPWR _03646_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_63_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07281_ data_array.data0\[8\]\[49\] net1389 net1295 data_array.data0\[11\]\[49\]
+ _04536_ VGND VGND VPWR VPWR _04537_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_100_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_151_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_151_clk
+ sky130_fd_sc_hd__clkbuf_8
X_09020_ net1987 net946 net418 VGND VGND VPWR VPWR _00775_ sky130_fd_sc_hd__mux2_1
X_06232_ tag_array.tag0\[8\]\[4\] net1373 net1279 tag_array.tag0\[11\]\[4\] _03582_
+ VGND VGND VPWR VPWR _03583_ sky130_fd_sc_hd__a221o_1
XFILLER_145_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06163_ tag_array.valid0\[1\] net1597 net1501 tag_array.valid0\[2\] VGND VGND VPWR
+ VPWR _03520_ sky130_fd_sc_hd__a22o_1
Xhold202 tag_array.tag1\[2\]\[12\] VGND VGND VPWR VPWR net1853 sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 data_array.data1\[1\]\[48\] VGND VGND VPWR VPWR net1864 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold224 data_array.data1\[2\]\[20\] VGND VGND VPWR VPWR net1875 sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 data_array.data0\[1\]\[53\] VGND VGND VPWR VPWR net1886 sky130_fd_sc_hd__dlygate4sd3_1
X_06094_ data_array.rdata0\[9\] net1139 net1114 data_array.rdata1\[9\] VGND VGND VPWR
+ VPWR net326 sky130_fd_sc_hd__a22o_1
Xhold246 data_array.data1\[0\]\[1\] VGND VGND VPWR VPWR net1897 sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 data_array.data0\[0\]\[29\] VGND VGND VPWR VPWR net1908 sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 data_array.data1\[2\]\[40\] VGND VGND VPWR VPWR net1919 sky130_fd_sc_hd__dlygate4sd3_1
Xhold279 data_array.data0\[4\]\[52\] VGND VGND VPWR VPWR net1930 sky130_fd_sc_hd__dlygate4sd3_1
X_09922_ net720 net3956 net602 VGND VGND VPWR VPWR _01672_ sky130_fd_sc_hd__mux2_1
Xfanout704 net705 VGND VGND VPWR VPWR net704 sky130_fd_sc_hd__clkbuf_2
Xfanout715 net717 VGND VGND VPWR VPWR net715 sky130_fd_sc_hd__buf_1
Xfanout726 net727 VGND VGND VPWR VPWR net726 sky130_fd_sc_hd__clkbuf_2
X_09853_ net1058 net3539 net380 VGND VGND VPWR VPWR _01603_ sky130_fd_sc_hd__mux2_1
Xfanout737 _05393_ VGND VGND VPWR VPWR net737 sky130_fd_sc_hd__clkbuf_2
Xfanout748 _05387_ VGND VGND VPWR VPWR net748 sky130_fd_sc_hd__clkbuf_2
XFILLER_113_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout759 _05381_ VGND VGND VPWR VPWR net759 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_146_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08804_ net3191 net1029 net448 VGND VGND VPWR VPWR _00562_ sky130_fd_sc_hd__mux2_1
X_09784_ net1073 net2701 net391 VGND VGND VPWR VPWR _01535_ sky130_fd_sc_hd__mux2_1
X_06996_ data_array.data0\[5\]\[23\] net1556 net1460 data_array.data0\[6\]\[23\] VGND
+ VGND VPWR VPWR _04278_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_163_3490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08735_ net783 net2395 net456 VGND VGND VPWR VPWR _00494_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05947_ net130 net1155 _03424_ _03425_ VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_1_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_124_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08666_ net760 net2367 net501 VGND VGND VPWR VPWR _00425_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_124_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05878_ net105 net1155 _03378_ _03379_ VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__a22o_1
X_07617_ data_array.data1\[9\]\[16\] net1545 net1449 data_array.data1\[10\]\[16\]
+ VGND VGND VPWR VPWR _04842_ sky130_fd_sc_hd__a22o_1
XFILLER_92_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08597_ net734 net3394 net529 VGND VGND VPWR VPWR _00356_ sky130_fd_sc_hd__mux2_1
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07548_ net1630 _04773_ _04777_ net1204 VGND VGND VPWR VPWR _04780_ sky130_fd_sc_hd__a22o_1
X_07479_ data_array.data1\[8\]\[3\] net1344 net1250 data_array.data1\[11\]\[3\] _04716_
+ VGND VGND VPWR VPWR _04717_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_142_clk clknet_5_30__leaf_clk VGND VGND VPWR VPWR clknet_leaf_142_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09218_ net708 net2084 net631 VGND VGND VPWR VPWR _00972_ sky130_fd_sc_hd__mux2_1
XFILLER_182_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10490_ net986 net4094 net348 VGND VGND VPWR VPWR _02235_ sky130_fd_sc_hd__mux2_1
XFILLER_182_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09149_ net947 net4064 net566 VGND VGND VPWR VPWR _00903_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12160_ clknet_leaf_108_clk _00968_ VGND VGND VPWR VPWR tag_array.tag0\[13\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_150_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11111_ net1075 net4522 net549 VGND VGND VPWR VPWR _02854_ sky130_fd_sc_hd__mux2_1
X_12091_ clknet_leaf_216_clk _00899_ VGND VGND VPWR VPWR data_array.data1\[14\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_9_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold780 data_array.data1\[6\]\[34\] VGND VGND VPWR VPWR net2431 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold791 tag_array.dirty0\[2\] VGND VGND VPWR VPWR net2442 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_1050 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11042_ net2505 net1092 net333 VGND VGND VPWR VPWR _02785_ sky130_fd_sc_hd__mux2_1
XFILLER_89_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_183_3866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_3877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2170 data_array.data0\[7\]\[54\] VGND VGND VPWR VPWR net3821 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_92_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2181 data_array.data1\[7\]\[43\] VGND VGND VPWR VPWR net3832 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2192 data_array.data1\[6\]\[47\] VGND VGND VPWR VPWR net3843 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12993_ clknet_leaf_15_clk _01687_ VGND VGND VPWR VPWR data_array.data0\[3\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1480 data_array.data1\[7\]\[17\] VGND VGND VPWR VPWR net3131 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_55_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1491 tag_array.tag1\[15\]\[24\] VGND VGND VPWR VPWR net3142 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11944_ clknet_leaf_48_clk _00752_ VGND VGND VPWR VPWR data_array.data0\[4\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_11875_ clknet_leaf_206_clk _00683_ VGND VGND VPWR VPWR data_array.data0\[5\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_10826_ net2213 net925 net502 VGND VGND VPWR VPWR _02571_ sky130_fd_sc_hd__mux2_1
X_13614_ clknet_leaf_235_clk _02243_ VGND VGND VPWR VPWR data_array.data0\[9\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_45_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13545_ clknet_leaf_88_clk _02174_ VGND VGND VPWR VPWR data_array.data1\[0\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
X_10757_ net944 net3900 net490 VGND VGND VPWR VPWR _02502_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_133_clk clknet_5_31__leaf_clk VGND VGND VPWR VPWR clknet_leaf_133_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_158_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13476_ clknet_leaf_158_clk _02106_ VGND VGND VPWR VPWR tag_array.tag0\[15\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_10688_ net2004 net965 net484 VGND VGND VPWR VPWR _02433_ sky130_fd_sc_hd__mux2_1
XFILLER_145_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12427_ clknet_leaf_20_clk _01121_ VGND VGND VPWR VPWR data_array.data0\[14\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_173_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput307 net307 VGND VGND VPWR VPWR mem_wdata[4] sky130_fd_sc_hd__buf_2
X_12358_ clknet_leaf_122_clk _00034_ VGND VGND VPWR VPWR data_array.rdata0\[40\] sky130_fd_sc_hd__dfxtp_1
Xoutput318 net318 VGND VGND VPWR VPWR mem_wdata[5] sky130_fd_sc_hd__buf_2
X_11309_ net1056 net2387 net798 VGND VGND VPWR VPWR _03052_ sky130_fd_sc_hd__mux2_1
XFILLER_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12289_ clknet_leaf_103_clk _01047_ VGND VGND VPWR VPWR tag_array.tag1\[13\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_142_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14028_ clknet_leaf_69_clk _02657_ VGND VGND VPWR VPWR data_array.data1\[6\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_06850_ data_array.data0\[4\]\[10\] net1411 net1317 data_array.data0\[7\]\[10\] _04144_
+ VGND VGND VPWR VPWR _04145_ sky130_fd_sc_hd__a221o_1
XFILLER_49_971 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_05801_ _03178_ _03179_ _03198_ _03229_ VGND VGND VPWR VPWR _03318_ sky130_fd_sc_hd__or4_1
XFILLER_95_587 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_887 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06781_ data_array.data0\[9\]\[4\] net1585 net1489 data_array.data0\[10\]\[4\] VGND
+ VGND VPWR VPWR _04082_ sky130_fd_sc_hd__a22o_1
X_08520_ net821 net812 net854 _05583_ VGND VGND VPWR VPWR _05585_ sky130_fd_sc_hd__or4b_1
X_05732_ fsm.tag_out1\[12\] net11 VGND VGND VPWR VPWR _03249_ sky130_fd_sc_hd__and2b_1
XFILLER_36_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08451_ net153 net88 net1640 VGND VGND VPWR VPWR _05537_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05663_ net2 fsm.tag_out0\[3\] VGND VGND VPWR VPWR _03180_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_102_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07402_ data_array.data0\[12\]\[60\] net1411 net1317 data_array.data0\[15\]\[60\]
+ _04646_ VGND VGND VPWR VPWR _04647_ sky130_fd_sc_hd__a221o_1
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08382_ net128 net63 net1648 VGND VGND VPWR VPWR _05491_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_82_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07333_ data_array.data0\[1\]\[54\] net1549 net1453 data_array.data0\[2\]\[54\] VGND
+ VGND VPWR VPWR _04584_ sky130_fd_sc_hd__a22o_1
XFILLER_52_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_124_clk clknet_5_27__leaf_clk VGND VGND VPWR VPWR clknet_leaf_124_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_176_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07264_ _04520_ _04521_ VGND VGND VPWR VPWR _00041_ sky130_fd_sc_hd__or2_1
XFILLER_137_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09003_ net1786 net1013 net424 VGND VGND VPWR VPWR _00758_ sky130_fd_sc_hd__mux2_1
X_06215_ tag_array.tag0\[1\]\[2\] net1560 net1464 tag_array.tag0\[2\]\[2\] VGND VGND
+ VPWR VPWR _03568_ sky130_fd_sc_hd__a22o_1
X_07195_ data_array.data0\[0\]\[41\] net1337 net1243 data_array.data0\[3\]\[41\] _04458_
+ VGND VGND VPWR VPWR _04459_ sky130_fd_sc_hd__a221o_1
X_06146_ data_array.rdata0\[61\] net1137 net1118 data_array.rdata1\[61\] VGND VGND
+ VPWR VPWR net320 sky130_fd_sc_hd__a22o_1
XFILLER_105_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_148_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06077_ net1161 net21 fsm.tag_out1\[21\] net1132 VGND VGND VPWR VPWR _03502_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_6_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout501 _05601_ VGND VGND VPWR VPWR net501 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_165_3530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_3541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09905_ net789 net2895 net602 VGND VGND VPWR VPWR _01655_ sky130_fd_sc_hd__mux2_1
XFILLER_99_871 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout512 net513 VGND VGND VPWR VPWR net512 sky130_fd_sc_hd__buf_2
Xfanout523 net525 VGND VGND VPWR VPWR net523 sky130_fd_sc_hd__clkbuf_8
Xfanout534 _05598_ VGND VGND VPWR VPWR net534 sky130_fd_sc_hd__clkbuf_4
Xfanout545 net546 VGND VGND VPWR VPWR net545 sky130_fd_sc_hd__buf_4
Xfanout556 net560 VGND VGND VPWR VPWR net556 sky130_fd_sc_hd__clkbuf_8
X_09836_ net867 net2737 net388 VGND VGND VPWR VPWR _01587_ sky130_fd_sc_hd__mux2_1
Xfanout567 net572 VGND VGND VPWR VPWR net567 sky130_fd_sc_hd__buf_4
Xfanout578 net581 VGND VGND VPWR VPWR net578 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_161_3449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout589 net590 VGND VGND VPWR VPWR net589 sky130_fd_sc_hd__buf_4
X_09767_ net2331 net718 net666 VGND VGND VPWR VPWR _01519_ sky130_fd_sc_hd__mux2_1
X_06979_ data_array.data0\[9\]\[22\] net1532 net1436 data_array.data0\[10\]\[22\]
+ VGND VGND VPWR VPWR _04262_ sky130_fd_sc_hd__a22o_1
XFILLER_26_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08718_ net3240 net750 net476 VGND VGND VPWR VPWR _00477_ sky130_fd_sc_hd__mux2_1
X_09698_ net696 net3916 net608 VGND VGND VPWR VPWR _01450_ sky130_fd_sc_hd__mux2_1
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_5_2__f_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_5_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_08649_ net1759 net728 net510 VGND VGND VPWR VPWR _00408_ sky130_fd_sc_hd__mux2_1
XFILLER_109_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11660_ clknet_leaf_99_clk _00468_ VGND VGND VPWR VPWR tag_array.tag1\[1\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_41_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10611_ net2203 net1016 net469 VGND VGND VPWR VPWR _02356_ sky130_fd_sc_hd__mux2_1
XFILLER_168_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11591_ clknet_leaf_132_clk _00399_ VGND VGND VPWR VPWR tag_array.tag1\[4\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_115_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_115_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13330_ clknet_leaf_235_clk _01960_ VGND VGND VPWR VPWR data_array.data0\[10\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
X_10542_ net1039 net3860 net455 VGND VGND VPWR VPWR _02287_ sky130_fd_sc_hd__mux2_1
XFILLER_183_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13261_ clknet_leaf_11_clk _01891_ VGND VGND VPWR VPWR data_array.data0\[11\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_137_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10473_ net1053 net4051 net348 VGND VGND VPWR VPWR _02218_ sky130_fd_sc_hd__mux2_1
XFILLER_109_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12212_ clknet_leaf_148_clk _00141_ VGND VGND VPWR VPWR fsm.tag_out0\[19\] sky130_fd_sc_hd__dfxtp_1
X_13192_ clknet_leaf_52_clk _00085_ VGND VGND VPWR VPWR data_array.rdata1\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12143_ clknet_leaf_159_clk _00951_ VGND VGND VPWR VPWR tag_array.tag0\[13\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_124_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12074_ clknet_leaf_122_clk _00882_ VGND VGND VPWR VPWR data_array.data1\[14\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_111_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11025_ net2376 net903 net338 VGND VGND VPWR VPWR _02769_ sky130_fd_sc_hd__mux2_1
XFILLER_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_86_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12976_ clknet_leaf_152_clk _01670_ VGND VGND VPWR VPWR tag_array.tag0\[4\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_45_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11927_ clknet_leaf_262_clk _00735_ VGND VGND VPWR VPWR data_array.data0\[4\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11858_ clknet_leaf_110_clk _00666_ VGND VGND VPWR VPWR data_array.data0\[7\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_19 _03480_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_106_clk clknet_5_25__leaf_clk VGND VGND VPWR VPWR clknet_leaf_106_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10809_ net1815 net994 net507 VGND VGND VPWR VPWR _02554_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11789_ clknet_leaf_13_clk _00597_ VGND VGND VPWR VPWR data_array.data0\[8\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_60_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13528_ clknet_leaf_267_clk _02157_ VGND VGND VPWR VPWR data_array.data1\[0\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_118_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13459_ clknet_leaf_164_clk _02089_ VGND VGND VPWR VPWR tag_array.tag0\[1\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_06000_ data_array.rdata1\[56\] net835 net844 VGND VGND VPWR VPWR _03461_ sky130_fd_sc_hd__a21o_1
XFILLER_141_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07951_ data_array.data1\[13\]\[46\] net1523 net1427 data_array.data1\[14\]\[46\]
+ VGND VGND VPWR VPWR _05146_ sky130_fd_sc_hd__a22o_1
XFILLER_99_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2906 data_array.data1\[6\]\[14\] VGND VGND VPWR VPWR net4557 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2917 data_array.data0\[9\]\[19\] VGND VGND VPWR VPWR net4568 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2928 data_array.data1\[9\]\[42\] VGND VGND VPWR VPWR net4579 sky130_fd_sc_hd__dlygate4sd3_1
X_06902_ data_array.data0\[9\]\[15\] net1584 net1488 data_array.data0\[10\]\[15\]
+ VGND VGND VPWR VPWR _04192_ sky130_fd_sc_hd__a22o_1
Xhold2939 tag_array.tag0\[1\]\[6\] VGND VGND VPWR VPWR net4590 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_143_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07882_ data_array.data1\[12\]\[40\] net1415 net1321 data_array.data1\[15\]\[40\]
+ _05082_ VGND VGND VPWR VPWR _05083_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_143_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09621_ net867 net2647 net396 VGND VGND VPWR VPWR _01373_ sky130_fd_sc_hd__mux2_1
X_06833_ net1194 _04123_ _04127_ net1620 VGND VGND VPWR VPWR _04130_ sky130_fd_sc_hd__a22o_1
XFILLER_28_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09552_ net720 net2830 net620 VGND VGND VPWR VPWR _01305_ sky130_fd_sc_hd__mux2_1
X_06764_ data_array.data0\[8\]\[2\] net1338 net1244 data_array.data0\[11\]\[2\] _04066_
+ VGND VGND VPWR VPWR _04067_ sky130_fd_sc_hd__a221o_1
X_08503_ net823 _05361_ VGND VGND VPWR VPWR _05572_ sky130_fd_sc_hd__or2_1
XFILLER_102_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05715_ _03173_ _03189_ _03190_ _03205_ VGND VGND VPWR VPWR _03232_ sky130_fd_sc_hd__or4_1
XFILLER_24_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09483_ net695 net3796 net653 VGND VGND VPWR VPWR _01236_ sky130_fd_sc_hd__mux2_1
X_06695_ tag_array.tag1\[5\]\[21\] net1592 net1496 tag_array.tag1\[6\]\[21\] VGND
+ VGND VPWR VPWR _04004_ sky130_fd_sc_hd__a22o_1
XFILLER_36_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08434_ net1123 _05525_ VGND VGND VPWR VPWR _05526_ sky130_fd_sc_hd__and2_1
XFILLER_51_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05646_ net24 fsm.tag_out0\[23\] VGND VGND VPWR VPWR _03163_ sky130_fd_sc_hd__xor2_1
XFILLER_168_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08365_ net1127 _05479_ VGND VGND VPWR VPWR _05480_ sky130_fd_sc_hd__and2_1
XFILLER_149_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07316_ data_array.data0\[0\]\[52\] net1357 net1263 data_array.data0\[3\]\[52\] _04568_
+ VGND VGND VPWR VPWR _04569_ sky130_fd_sc_hd__a221o_1
X_08296_ net1129 _05433_ VGND VGND VPWR VPWR _05434_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_119_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07247_ data_array.data0\[13\]\[46\] net1532 net1436 data_array.data0\[14\]\[46\]
+ VGND VGND VPWR VPWR _04506_ sky130_fd_sc_hd__a22o_1
XFILLER_165_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_2_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_2_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_139_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07178_ data_array.data0\[12\]\[40\] net1413 net1319 data_array.data0\[15\]\[40\]
+ _04442_ VGND VGND VPWR VPWR _04443_ sky130_fd_sc_hd__a221o_1
XFILLER_105_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06129_ data_array.rdata0\[44\] net1139 net1115 data_array.rdata1\[44\] VGND VGND
+ VPWR VPWR net301 sky130_fd_sc_hd__a22o_1
XFILLER_105_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1307 net1309 VGND VGND VPWR VPWR net1307 sky130_fd_sc_hd__clkbuf_4
Xfanout1318 net1319 VGND VGND VPWR VPWR net1318 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_180_3814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1329 net1331 VGND VGND VPWR VPWR net1329 sky130_fd_sc_hd__clkbuf_4
Xfanout331 net332 VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_180_3825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout342 net343 VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__buf_4
Xfanout353 _03130_ VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__buf_1
Xfanout364 net365 VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__buf_4
Xfanout375 net376 VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__buf_4
Xfanout386 net387 VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__clkbuf_8
X_09819_ net933 net2893 net392 VGND VGND VPWR VPWR _01570_ sky130_fd_sc_hd__mux2_1
Xfanout397 net401 VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__buf_4
XFILLER_98_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12830_ clknet_leaf_129_clk _01524_ VGND VGND VPWR VPWR tag_array.tag1\[0\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_98_1059 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12761_ clknet_leaf_177_clk _01455_ VGND VGND VPWR VPWR tag_array.tag0\[6\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_6_Left_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_178_3776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ clknet_leaf_177_clk _03121_ VGND VGND VPWR VPWR lru_array.lru_mem\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_178_3787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ clknet_leaf_171_clk _00520_ VGND VGND VPWR VPWR tag_array.tag0\[9\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_43_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12692_ clknet_leaf_107_clk _01386_ VGND VGND VPWR VPWR tag_array.tag0\[8\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_42_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14431_ clknet_leaf_66_clk _03054_ VGND VGND VPWR VPWR data_array.data1\[7\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_11643_ clknet_leaf_127_clk _00451_ VGND VGND VPWR VPWR tag_array.tag1\[2\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14362_ clknet_leaf_84_clk _02985_ VGND VGND VPWR VPWR data_array.data1\[10\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_11574_ clknet_leaf_99_clk _00382_ VGND VGND VPWR VPWR tag_array.tag1\[5\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput17 cpu_addr[24] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_2
XFILLER_168_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput28 cpu_addr[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_4
X_10525_ net1107 net4549 net453 VGND VGND VPWR VPWR _02270_ sky130_fd_sc_hd__mux2_1
X_13313_ clknet_leaf_22_clk _01943_ VGND VGND VPWR VPWR data_array.data0\[10\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput39 cpu_wdata[14] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_1
X_14293_ clknet_leaf_199_clk _02922_ VGND VGND VPWR VPWR data_array.data1\[11\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13244_ clknet_leaf_249_clk _01874_ VGND VGND VPWR VPWR data_array.data0\[11\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_10456_ net1964 net353 net467 VGND VGND VPWR VPWR _02202_ sky130_fd_sc_hd__mux2_1
XFILLER_109_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13175_ clknet_leaf_81_clk _00067_ VGND VGND VPWR VPWR data_array.rdata1\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_151_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10387_ net1897 net1104 net661 VGND VGND VPWR VPWR _02133_ sky130_fd_sc_hd__mux2_1
X_12126_ clknet_leaf_145_clk _00934_ VGND VGND VPWR VPWR tag_array.tag0\[12\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_97_627 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12057_ clknet_leaf_36_clk _00865_ VGND VGND VPWR VPWR data_array.data1\[14\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_77_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11008_ net2555 net971 net336 VGND VGND VPWR VPWR _02752_ sky130_fd_sc_hd__mux2_1
XFILLER_77_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12959_ clknet_leaf_225_clk _01653_ VGND VGND VPWR VPWR data_array.data0\[13\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_93_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06480_ tag_array.tag1\[0\]\[1\] net1401 net1307 tag_array.tag1\[3\]\[1\] _03808_
+ VGND VGND VPWR VPWR _03809_ sky130_fd_sc_hd__a221o_1
XFILLER_33_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08150_ tag_array.dirty1\[8\] net1350 net1256 tag_array.dirty1\[11\] _05326_ VGND
+ VGND VPWR VPWR _05327_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_99_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07101_ data_array.data0\[12\]\[33\] net1396 net1302 data_array.data0\[15\]\[33\]
+ _04372_ VGND VGND VPWR VPWR _04373_ sky130_fd_sc_hd__a221o_1
XFILLER_119_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08081_ data_array.data1\[5\]\[58\] net1550 net1454 data_array.data1\[6\]\[58\] VGND
+ VGND VPWR VPWR _05264_ sky130_fd_sc_hd__a22o_1
Xclkload200 clknet_leaf_163_clk VGND VGND VPWR VPWR clkload200/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload211 clknet_leaf_119_clk VGND VGND VPWR VPWR clkload211/X sky130_fd_sc_hd__clkbuf_4
XFILLER_146_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload222 clknet_leaf_159_clk VGND VGND VPWR VPWR clkload222/Y sky130_fd_sc_hd__bufinv_16
Xclkload233 clknet_leaf_131_clk VGND VGND VPWR VPWR clkload233/Y sky130_fd_sc_hd__inv_16
XFILLER_162_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07032_ net1167 _04305_ _04309_ net1214 VGND VGND VPWR VPWR _04311_ sky130_fd_sc_hd__a22o_1
Xclkload244 clknet_leaf_141_clk VGND VGND VPWR VPWR clkload244/Y sky130_fd_sc_hd__clkinv_2
XFILLER_173_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2703 data_array.data0\[15\]\[44\] VGND VGND VPWR VPWR net4354 sky130_fd_sc_hd__dlygate4sd3_1
X_08983_ net3018 net1093 net423 VGND VGND VPWR VPWR _00738_ sky130_fd_sc_hd__mux2_1
Xhold2714 data_array.data0\[14\]\[14\] VGND VGND VPWR VPWR net4365 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_110_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2725 data_array.data1\[15\]\[8\] VGND VGND VPWR VPWR net4376 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07934_ net1227 _05125_ _05129_ net1180 VGND VGND VPWR VPWR _05131_ sky130_fd_sc_hd__a22o_1
Xhold2736 tag_array.tag1\[14\]\[11\] VGND VGND VPWR VPWR net4387 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2747 tag_array.tag1\[9\]\[20\] VGND VGND VPWR VPWR net4398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2758 data_array.data1\[11\]\[42\] VGND VGND VPWR VPWR net4409 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2769 data_array.data1\[3\]\[6\] VGND VGND VPWR VPWR net4420 sky130_fd_sc_hd__dlygate4sd3_1
X_07865_ data_array.data1\[5\]\[38\] net1588 net1492 data_array.data1\[6\]\[38\] VGND
+ VGND VPWR VPWR _05068_ sky130_fd_sc_hd__a22o_1
XFILLER_29_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09604_ net933 net4354 net400 VGND VGND VPWR VPWR _01356_ sky130_fd_sc_hd__mux2_1
XFILLER_28_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06816_ data_array.data0\[1\]\[7\] net1601 net1505 data_array.data0\[2\]\[7\] VGND
+ VGND VPWR VPWR _04114_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_27_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07796_ data_array.data1\[0\]\[32\] net1330 net1236 data_array.data1\[3\]\[32\] _05004_
+ VGND VGND VPWR VPWR _05005_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_27_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06747_ _04050_ _04051_ VGND VGND VPWR VPWR _00000_ sky130_fd_sc_hd__or2_2
X_09535_ net789 net3251 net618 VGND VGND VPWR VPWR _01288_ sky130_fd_sc_hd__mux2_1
X_09466_ net765 net3695 net658 VGND VGND VPWR VPWR _01219_ sky130_fd_sc_hd__mux2_1
X_06678_ tag_array.tag1\[0\]\[19\] net1404 net1310 tag_array.tag1\[3\]\[19\] _03988_
+ VGND VGND VPWR VPWR _03989_ sky130_fd_sc_hd__a221o_1
XFILLER_40_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_3359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05629_ net4624 _03148_ net229 VGND VGND VPWR VPWR _00186_ sky130_fd_sc_hd__a21o_1
X_08417_ net1834 net921 net691 VGND VGND VPWR VPWR _00268_ sky130_fd_sc_hd__mux2_1
XFILLER_12_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09397_ net1079 net2483 net580 VGND VGND VPWR VPWR _01150_ sky130_fd_sc_hd__mux2_1
X_08348_ net2089 net1013 net693 VGND VGND VPWR VPWR _00245_ sky130_fd_sc_hd__mux2_1
XFILLER_132_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08279_ net1931 net1105 net686 VGND VGND VPWR VPWR _00222_ sky130_fd_sc_hd__mux2_1
XFILLER_22_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10310_ net2294 net922 net641 VGND VGND VPWR VPWR _02057_ sky130_fd_sc_hd__mux2_1
XFILLER_138_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11290_ net871 net2401 net683 VGND VGND VPWR VPWR _03033_ sky130_fd_sc_hd__mux2_1
XFILLER_152_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10241_ net780 net2779 net595 VGND VGND VPWR VPWR _01988_ sky130_fd_sc_hd__mux2_1
XFILLER_121_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10172_ net856 net2804 net364 VGND VGND VPWR VPWR _01920_ sky130_fd_sc_hd__mux2_1
Xfanout1104 net1107 VGND VGND VPWR VPWR net1104 sky130_fd_sc_hd__clkbuf_2
Xfanout1115 net1116 VGND VGND VPWR VPWR net1115 sky130_fd_sc_hd__buf_4
Xfanout1126 net1130 VGND VGND VPWR VPWR net1126 sky130_fd_sc_hd__clkbuf_2
Xfanout1137 net1138 VGND VGND VPWR VPWR net1137 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1148 net1149 VGND VGND VPWR VPWR net1148 sky130_fd_sc_hd__buf_4
Xfanout1159 net1160 VGND VGND VPWR VPWR net1159 sky130_fd_sc_hd__clkbuf_2
XFILLER_102_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_362 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13931_ clknet_leaf_256_clk _02560_ VGND VGND VPWR VPWR data_array.data1\[4\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_822 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13862_ clknet_leaf_69_clk _02491_ VGND VGND VPWR VPWR data_array.data1\[3\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_170_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12813_ clknet_leaf_195_clk _01507_ VGND VGND VPWR VPWR tag_array.tag1\[0\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_13793_ clknet_leaf_267_clk _02422_ VGND VGND VPWR VPWR data_array.data1\[2\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12744_ clknet_leaf_155_clk _01438_ VGND VGND VPWR VPWR tag_array.tag0\[5\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_179_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12675_ clknet_leaf_234_clk _01369_ VGND VGND VPWR VPWR data_array.data0\[15\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_147_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14414_ clknet_leaf_179_clk _03037_ VGND VGND VPWR VPWR lru_array.lru_mem\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_169_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11626_ clknet_leaf_128_clk _00434_ VGND VGND VPWR VPWR tag_array.tag1\[3\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_156_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14345_ clknet_leaf_184_clk _00187_ _00190_ VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__dfrtp_1
X_11557_ clknet_leaf_129_clk _00365_ VGND VGND VPWR VPWR tag_array.tag1\[6\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold609 data_array.data0\[8\]\[28\] VGND VGND VPWR VPWR net2260 sky130_fd_sc_hd__dlygate4sd3_1
X_10508_ net913 net2488 net349 VGND VGND VPWR VPWR _02253_ sky130_fd_sc_hd__mux2_1
X_14276_ clknet_leaf_119_clk _02905_ VGND VGND VPWR VPWR data_array.data1\[12\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
X_11488_ clknet_leaf_153_clk _00297_ VGND VGND VPWR VPWR tag_array.valid0\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_109_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10439_ net2663 net898 net661 VGND VGND VPWR VPWR _02185_ sky130_fd_sc_hd__mux2_1
X_13227_ clknet_leaf_227_clk _01857_ VGND VGND VPWR VPWR data_array.data0\[11\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_171_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13158_ clknet_leaf_232_clk _01852_ VGND VGND VPWR VPWR tag_array.tag1\[8\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_98_958 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ clknet_leaf_21_clk _00917_ VGND VGND VPWR VPWR data_array.data1\[14\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_72_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13089_ clknet_leaf_121_clk _01783_ VGND VGND VPWR VPWR data_array.data1\[13\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
X_05980_ net142 net1155 _03446_ _03447_ VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__a22o_1
Xhold1309 tag_array.tag1\[15\]\[7\] VGND VGND VPWR VPWR net2960 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07650_ data_array.data1\[13\]\[19\] net1584 net1488 data_array.data1\[14\]\[19\]
+ VGND VGND VPWR VPWR _04872_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_69_Left_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06601_ tag_array.tag1\[0\]\[12\] net1401 net1307 tag_array.tag1\[3\]\[12\] _03918_
+ VGND VGND VPWR VPWR _03919_ sky130_fd_sc_hd__a221o_1
X_07581_ net1631 _04803_ _04807_ net1205 VGND VGND VPWR VPWR _04810_ sky130_fd_sc_hd__a22o_1
XFILLER_25_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09320_ net700 net3757 net552 VGND VGND VPWR VPWR _01074_ sky130_fd_sc_hd__mux2_1
X_06532_ tag_array.tag1\[9\]\[6\] net1552 net1456 tag_array.tag1\[10\]\[6\] VGND VGND
+ VPWR VPWR _03856_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_138_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09251_ net774 net2617 net570 VGND VGND VPWR VPWR _01005_ sky130_fd_sc_hd__mux2_1
XFILLER_21_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06463_ tag_array.tag1\[8\]\[0\] net1386 net1292 tag_array.tag1\[11\]\[0\] _03792_
+ VGND VGND VPWR VPWR _03793_ sky130_fd_sc_hd__a221o_1
X_08202_ net782 net4307 net797 VGND VGND VPWR VPWR _00198_ sky130_fd_sc_hd__mux2_1
XFILLER_21_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09182_ net753 net3785 net628 VGND VGND VPWR VPWR _00936_ sky130_fd_sc_hd__mux2_1
X_06394_ net1230 _03725_ _03729_ net1182 VGND VGND VPWR VPWR _03731_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_79_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08133_ _05310_ _05311_ VGND VGND VPWR VPWR _00122_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_32_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1052 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_78_Left_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_151_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08064_ data_array.data1\[0\]\[56\] net1340 net1246 data_array.data1\[3\]\[56\] _05248_
+ VGND VGND VPWR VPWR _05249_ sky130_fd_sc_hd__a221o_1
XFILLER_162_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07015_ data_array.data0\[0\]\[25\] net1329 net1235 data_array.data0\[3\]\[25\] _04294_
+ VGND VGND VPWR VPWR _04295_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_112_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1039 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2500 tag_array.tag1\[10\]\[20\] VGND VGND VPWR VPWR net4151 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2511 data_array.data0\[7\]\[35\] VGND VGND VPWR VPWR net4162 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2522 tag_array.tag1\[15\]\[5\] VGND VGND VPWR VPWR net4173 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2533 data_array.data0\[12\]\[38\] VGND VGND VPWR VPWR net4184 sky130_fd_sc_hd__dlygate4sd3_1
X_08966_ net902 net3125 net429 VGND VGND VPWR VPWR _00722_ sky130_fd_sc_hd__mux2_1
Xhold2544 data_array.data0\[7\]\[32\] VGND VGND VPWR VPWR net4195 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1810 data_array.data1\[9\]\[1\] VGND VGND VPWR VPWR net3461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2555 tag_array.tag1\[7\]\[3\] VGND VGND VPWR VPWR net4206 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2566 data_array.data1\[12\]\[15\] VGND VGND VPWR VPWR net4217 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1821 tag_array.tag0\[1\]\[24\] VGND VGND VPWR VPWR net3472 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_87_Left_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07917_ data_array.data1\[0\]\[43\] net1378 net1284 data_array.data1\[3\]\[43\] _05114_
+ VGND VGND VPWR VPWR _05115_ sky130_fd_sc_hd__a221o_1
Xhold2577 data_array.data0\[6\]\[3\] VGND VGND VPWR VPWR net4228 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1832 data_array.data0\[12\]\[24\] VGND VGND VPWR VPWR net3483 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2588 data_array.data1\[5\]\[1\] VGND VGND VPWR VPWR net4239 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1843 data_array.data1\[5\]\[26\] VGND VGND VPWR VPWR net3494 sky130_fd_sc_hd__dlygate4sd3_1
X_08897_ net917 net2519 net438 VGND VGND VPWR VPWR _00654_ sky130_fd_sc_hd__mux2_1
Xhold1854 tag_array.tag1\[8\]\[7\] VGND VGND VPWR VPWR net3505 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_95_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_95_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_29_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2599 tag_array.tag0\[9\]\[23\] VGND VGND VPWR VPWR net4250 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1865 tag_array.tag0\[6\]\[17\] VGND VGND VPWR VPWR net3516 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1876 data_array.data0\[7\]\[62\] VGND VGND VPWR VPWR net3527 sky130_fd_sc_hd__dlygate4sd3_1
X_07848_ data_array.data1\[9\]\[37\] net1544 net1448 data_array.data1\[10\]\[37\]
+ VGND VGND VPWR VPWR _05052_ sky130_fd_sc_hd__a22o_1
Xhold1887 tag_array.tag1\[13\]\[4\] VGND VGND VPWR VPWR net3538 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_162_Right_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1898 data_array.data1\[14\]\[23\] VGND VGND VPWR VPWR net3549 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07779_ net1630 _04983_ _04987_ net1204 VGND VGND VPWR VPWR _04990_ sky130_fd_sc_hd__a22o_1
X_09518_ net755 net2098 net622 VGND VGND VPWR VPWR _01271_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_175_3724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10790_ net2068 net1071 net510 VGND VGND VPWR VPWR _02535_ sky130_fd_sc_hd__mux2_1
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09449_ net871 net2794 net588 VGND VGND VPWR VPWR _01202_ sky130_fd_sc_hd__mux2_1
XFILLER_24_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_96_Left_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12460_ clknet_leaf_84_clk _01154_ VGND VGND VPWR VPWR data_array.data1\[9\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11411_ clknet_leaf_230_clk _00221_ VGND VGND VPWR VPWR data_array.data0\[0\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_138_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12391_ clknet_leaf_61_clk _01085_ VGND VGND VPWR VPWR data_array.data0\[14\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_153_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11342_ net925 net4444 net795 VGND VGND VPWR VPWR _03085_ sky130_fd_sc_hd__mux2_1
X_14130_ clknet_leaf_93_clk _02759_ VGND VGND VPWR VPWR data_array.data0\[1\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_181_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14061_ clknet_leaf_215_clk _02690_ VGND VGND VPWR VPWR data_array.data1\[6\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
X_11273_ net937 net4231 net680 VGND VGND VPWR VPWR _03016_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13012_ clknet_leaf_238_clk _01706_ VGND VGND VPWR VPWR data_array.data0\[3\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_10224_ net910 net4088 net361 VGND VGND VPWR VPWR _01971_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10155_ net927 net3052 net362 VGND VGND VPWR VPWR _01903_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_468 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10086_ net2300 net779 _05557_ VGND VGND VPWR VPWR _01835_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_86_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_86_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_48_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13914_ clknet_leaf_18_clk _02543_ VGND VGND VPWR VPWR data_array.data1\[4\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13845_ clknet_leaf_200_clk _02474_ VGND VGND VPWR VPWR data_array.data1\[3\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_774 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13776_ clknet_leaf_19_clk _02405_ VGND VGND VPWR VPWR data_array.data1\[2\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_10988_ net1850 net1048 net341 VGND VGND VPWR VPWR _02732_ sky130_fd_sc_hd__mux2_1
X_12727_ clknet_leaf_169_clk _01421_ VGND VGND VPWR VPWR tag_array.tag0\[7\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_175_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12658_ clknet_leaf_124_clk _01352_ VGND VGND VPWR VPWR data_array.data0\[15\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_96_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11609_ clknet_leaf_97_clk _00417_ VGND VGND VPWR VPWR tag_array.tag1\[3\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_157_974 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12589_ clknet_leaf_155_clk _01283_ VGND VGND VPWR VPWR tag_array.tag0\[10\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_10_clk clknet_5_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_8
X_14328_ clknet_leaf_75_clk _02957_ VGND VGND VPWR VPWR data_array.data1\[11\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold406 data_array.data0\[1\]\[17\] VGND VGND VPWR VPWR net2057 sky130_fd_sc_hd__dlygate4sd3_1
Xhold417 data_array.data1\[4\]\[10\] VGND VGND VPWR VPWR net2068 sky130_fd_sc_hd__dlygate4sd3_1
Xhold428 data_array.data0\[8\]\[56\] VGND VGND VPWR VPWR net2079 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold439 data_array.data1\[15\]\[13\] VGND VGND VPWR VPWR net2090 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14259_ clknet_leaf_43_clk _02888_ VGND VGND VPWR VPWR data_array.data1\[12\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout908 net911 VGND VGND VPWR VPWR net908 sky130_fd_sc_hd__clkbuf_2
XFILLER_124_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout919 _05516_ VGND VGND VPWR VPWR net919 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_70_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08820_ net2264 net965 net448 VGND VGND VPWR VPWR _00578_ sky130_fd_sc_hd__mux2_1
XFILLER_97_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1106 tag_array.tag0\[7\]\[12\] VGND VGND VPWR VPWR net2757 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1117 data_array.data0\[10\]\[36\] VGND VGND VPWR VPWR net2768 sky130_fd_sc_hd__dlygate4sd3_1
X_05963_ data_array.rdata0\[44\] net852 net1148 VGND VGND VPWR VPWR _03436_ sky130_fd_sc_hd__o21a_1
Xhold1128 tag_array.tag0\[2\]\[3\] VGND VGND VPWR VPWR net2779 sky130_fd_sc_hd__dlygate4sd3_1
X_08751_ net718 net2343 net458 VGND VGND VPWR VPWR _00510_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_77_clk clknet_5_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_77_clk sky130_fd_sc_hd__clkbuf_8
Xhold1139 data_array.data1\[2\]\[41\] VGND VGND VPWR VPWR net2790 sky130_fd_sc_hd__dlygate4sd3_1
X_07702_ net1196 _04913_ _04917_ net1622 VGND VGND VPWR VPWR _04920_ sky130_fd_sc_hd__a22o_1
Xfanout1490 net1491 VGND VGND VPWR VPWR net1490 sky130_fd_sc_hd__clkbuf_4
X_05894_ data_array.rdata0\[21\] net848 net1144 VGND VGND VPWR VPWR _03390_ sky130_fd_sc_hd__o21a_1
XFILLER_39_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08682_ net695 net2184 net494 VGND VGND VPWR VPWR _00441_ sky130_fd_sc_hd__mux2_1
XFILLER_81_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07633_ data_array.data1\[8\]\[17\] net1336 net1242 data_array.data1\[11\]\[17\]
+ _04856_ VGND VGND VPWR VPWR _04857_ sky130_fd_sc_hd__a221o_1
XFILLER_54_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07564_ data_array.data1\[1\]\[11\] net1576 net1480 data_array.data1\[2\]\[11\] VGND
+ VGND VPWR VPWR _04794_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_105_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_105_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_532 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06515_ net1220 _03835_ _03839_ net1174 VGND VGND VPWR VPWR _03841_ sky130_fd_sc_hd__a22o_1
X_09303_ net766 net2867 net546 VGND VGND VPWR VPWR _01057_ sky130_fd_sc_hd__mux2_1
X_07495_ _04730_ _04731_ VGND VGND VPWR VPWR _00108_ sky130_fd_sc_hd__or2_1
XFILLER_22_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09234_ net744 net3665 net645 VGND VGND VPWR VPWR _00988_ sky130_fd_sc_hd__mux2_1
X_06446_ tag_array.tag0\[5\]\[23\] net1602 net1506 tag_array.tag0\[6\]\[23\] VGND
+ VGND VPWR VPWR _03778_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_170_3621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09165_ net882 net4374 net567 VGND VGND VPWR VPWR _00919_ sky130_fd_sc_hd__mux2_1
XFILLER_21_298 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06377_ tag_array.tag0\[4\]\[17\] net1412 net1318 tag_array.tag0\[7\]\[17\] _03714_
+ VGND VGND VPWR VPWR _03715_ sky130_fd_sc_hd__a221o_1
XFILLER_119_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08116_ data_array.data1\[9\]\[61\] net1545 net1449 data_array.data1\[10\]\[61\]
+ VGND VGND VPWR VPWR _05296_ sky130_fd_sc_hd__a22o_1
XFILLER_147_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09096_ net902 net2780 net413 VGND VGND VPWR VPWR _00850_ sky130_fd_sc_hd__mux2_1
XFILLER_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08047_ data_array.data1\[12\]\[55\] net1344 net1250 data_array.data1\[15\]\[55\]
+ _05232_ VGND VGND VPWR VPWR _05233_ sky130_fd_sc_hd__a221o_1
XFILLER_79_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold940 data_array.data0\[11\]\[17\] VGND VGND VPWR VPWR net2591 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold951 data_array.data0\[13\]\[48\] VGND VGND VPWR VPWR net2602 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold962 tag_array.tag1\[5\]\[10\] VGND VGND VPWR VPWR net2613 sky130_fd_sc_hd__dlygate4sd3_1
Xhold973 data_array.data0\[4\]\[58\] VGND VGND VPWR VPWR net2624 sky130_fd_sc_hd__dlygate4sd3_1
Xhold984 tag_array.dirty1\[14\] VGND VGND VPWR VPWR net2635 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_168_3583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold995 tag_array.tag0\[2\]\[17\] VGND VGND VPWR VPWR net2646 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_168_3594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09998_ net1095 net2773 net562 VGND VGND VPWR VPWR _01747_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2330 data_array.data0\[15\]\[59\] VGND VGND VPWR VPWR net3981 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2341 data_array.data1\[2\]\[55\] VGND VGND VPWR VPWR net3992 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2352 data_array.data1\[12\]\[22\] VGND VGND VPWR VPWR net4003 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08949_ net970 net2323 net426 VGND VGND VPWR VPWR _00705_ sky130_fd_sc_hd__mux2_1
Xhold2363 data_array.data1\[11\]\[55\] VGND VGND VPWR VPWR net4014 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_68_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_68_clk sky130_fd_sc_hd__clkbuf_8
Xhold2374 data_array.data0\[3\]\[6\] VGND VGND VPWR VPWR net4025 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2385 data_array.data0\[12\]\[27\] VGND VGND VPWR VPWR net4036 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1640 tag_array.tag1\[13\]\[1\] VGND VGND VPWR VPWR net3291 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2396 data_array.data0\[13\]\[17\] VGND VGND VPWR VPWR net4047 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1651 data_array.data0\[6\]\[40\] VGND VGND VPWR VPWR net3302 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1662 data_array.data1\[14\]\[40\] VGND VGND VPWR VPWR net3313 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11960_ clknet_leaf_11_clk _00768_ VGND VGND VPWR VPWR data_array.data0\[4\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1673 data_array.data1\[13\]\[5\] VGND VGND VPWR VPWR net3324 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1684 tag_array.tag1\[14\]\[16\] VGND VGND VPWR VPWR net3335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1695 data_array.data1\[10\]\[20\] VGND VGND VPWR VPWR net3346 sky130_fd_sc_hd__dlygate4sd3_1
X_10911_ net1098 net4126 net531 VGND VGND VPWR VPWR _02656_ sky130_fd_sc_hd__mux2_1
XFILLER_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11891_ clknet_leaf_52_clk _00699_ VGND VGND VPWR VPWR data_array.data0\[5\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_13630_ clknet_leaf_13_clk _02259_ VGND VGND VPWR VPWR data_array.data0\[9\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
X_10842_ net2104 net862 net510 VGND VGND VPWR VPWR _02587_ sky130_fd_sc_hd__mux2_1
XFILLER_44_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13561_ clknet_leaf_202_clk _02190_ VGND VGND VPWR VPWR data_array.data1\[0\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
X_10773_ net883 net3148 net491 VGND VGND VPWR VPWR _02518_ sky130_fd_sc_hd__mux2_1
XFILLER_12_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12512_ clknet_leaf_178_clk _01206_ VGND VGND VPWR VPWR lru_array.lru_mem\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_157_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13492_ clknet_leaf_159_clk _02122_ VGND VGND VPWR VPWR tag_array.tag0\[15\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_157_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12443_ clknet_leaf_205_clk _01137_ VGND VGND VPWR VPWR data_array.data0\[14\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_139_985 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12374_ clknet_leaf_12_clk _00051_ VGND VGND VPWR VPWR data_array.rdata0\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_165_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14113_ clknet_leaf_0_clk _02742_ VGND VGND VPWR VPWR data_array.data0\[1\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_158_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11325_ net994 net4358 net800 VGND VGND VPWR VPWR _03068_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14044_ clknet_leaf_123_clk _02673_ VGND VGND VPWR VPWR data_array.data1\[6\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_158_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11256_ net1005 net4050 net674 VGND VGND VPWR VPWR _02999_ sky130_fd_sc_hd__mux2_1
X_10207_ net977 net4236 net359 VGND VGND VPWR VPWR _01954_ sky130_fd_sc_hd__mux2_1
X_11187_ net1025 net4186 net652 VGND VGND VPWR VPWR _02930_ sky130_fd_sc_hd__mux2_1
X_10138_ net993 net4285 net367 VGND VGND VPWR VPWR _01886_ sky130_fd_sc_hd__mux2_1
XFILLER_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_59_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_59_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_89_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10069_ net748 net2909 net600 VGND VGND VPWR VPWR _01818_ sky130_fd_sc_hd__mux2_1
XFILLER_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_644 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13828_ clknet_leaf_115_clk _02457_ VGND VGND VPWR VPWR data_array.data1\[2\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13759_ clknet_leaf_17_clk _02388_ VGND VGND VPWR VPWR data_array.data1\[1\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06300_ tag_array.tag0\[4\]\[10\] net1405 net1311 tag_array.tag0\[7\]\[10\] _03644_
+ VGND VGND VPWR VPWR _03645_ sky130_fd_sc_hd__a221o_1
XFILLER_31_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07280_ data_array.data0\[9\]\[49\] net1580 net1484 data_array.data0\[10\]\[49\]
+ VGND VGND VPWR VPWR _04536_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_63_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1030 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06231_ tag_array.tag0\[9\]\[4\] net1564 net1468 tag_array.tag0\[10\]\[4\] VGND VGND
+ VPWR VPWR _03582_ sky130_fd_sc_hd__a22o_1
XFILLER_117_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06162_ net28 net29 VGND VGND VPWR VPWR _03519_ sky130_fd_sc_hd__or2_2
XFILLER_117_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold203 data_array.data0\[1\]\[40\] VGND VGND VPWR VPWR net1854 sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 data_array.data1\[8\]\[43\] VGND VGND VPWR VPWR net1865 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_160_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold225 data_array.data1\[4\]\[63\] VGND VGND VPWR VPWR net1876 sky130_fd_sc_hd__dlygate4sd3_1
X_06093_ data_array.rdata0\[8\] net1135 net1112 data_array.rdata1\[8\] VGND VGND VPWR
+ VPWR net325 sky130_fd_sc_hd__a22o_1
Xhold236 data_array.data1\[2\]\[58\] VGND VGND VPWR VPWR net1887 sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 data_array.data1\[1\]\[2\] VGND VGND VPWR VPWR net1898 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 data_array.data0\[2\]\[60\] VGND VGND VPWR VPWR net1909 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold269 tag_array.tag1\[0\]\[24\] VGND VGND VPWR VPWR net1920 sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ net722 net2812 net603 VGND VGND VPWR VPWR _01671_ sky130_fd_sc_hd__mux2_1
Xfanout705 _05409_ VGND VGND VPWR VPWR net705 sky130_fd_sc_hd__clkbuf_2
Xfanout716 net717 VGND VGND VPWR VPWR net716 sky130_fd_sc_hd__clkbuf_2
Xfanout727 _05397_ VGND VGND VPWR VPWR net727 sky130_fd_sc_hd__dlymetal6s2s_1
X_09852_ net1061 net2586 net384 VGND VGND VPWR VPWR _01602_ sky130_fd_sc_hd__mux2_1
Xfanout738 _05391_ VGND VGND VPWR VPWR net738 sky130_fd_sc_hd__clkbuf_2
Xfanout749 _05387_ VGND VGND VPWR VPWR net749 sky130_fd_sc_hd__buf_1
X_08803_ net1740 net1032 net447 VGND VGND VPWR VPWR _00561_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_146_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ net1079 net3687 net387 VGND VGND VPWR VPWR _01534_ sky130_fd_sc_hd__mux2_1
XFILLER_105_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1001 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06995_ data_array.data0\[8\]\[23\] net1371 net1277 data_array.data0\[11\]\[23\]
+ _04276_ VGND VGND VPWR VPWR _04277_ sky130_fd_sc_hd__a221o_1
XFILLER_39_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_163_3491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08734_ net786 net3063 net455 VGND VGND VPWR VPWR _00493_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05946_ data_array.rdata1\[38\] net832 net841 VGND VGND VPWR VPWR _03425_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_107_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08665_ net764 net3661 net500 VGND VGND VPWR VPWR _00424_ sky130_fd_sc_hd__mux2_1
X_05877_ data_array.rdata1\[15\] net832 net841 VGND VGND VPWR VPWR _03379_ sky130_fd_sc_hd__a21o_1
XFILLER_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_124_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07616_ _04840_ _04841_ VGND VGND VPWR VPWR _00070_ sky130_fd_sc_hd__or2_1
X_08596_ net740 net3940 net536 VGND VGND VPWR VPWR _00355_ sky130_fd_sc_hd__mux2_1
XFILLER_35_880 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07547_ data_array.data1\[0\]\[9\] net1389 net1295 data_array.data1\[3\]\[9\] _04778_
+ VGND VGND VPWR VPWR _04779_ sky130_fd_sc_hd__a221o_1
XFILLER_179_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07478_ data_array.data1\[9\]\[3\] net1535 net1439 data_array.data1\[10\]\[3\] VGND
+ VGND VPWR VPWR _04716_ sky130_fd_sc_hd__a22o_1
XFILLER_167_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09217_ net713 net2956 net630 VGND VGND VPWR VPWR _00971_ sky130_fd_sc_hd__mux2_1
X_06429_ tag_array.tag0\[9\]\[22\] net1565 net1469 tag_array.tag0\[10\]\[22\] VGND
+ VGND VPWR VPWR _03762_ sky130_fd_sc_hd__a22o_1
XFILLER_6_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09148_ net951 net3313 net576 VGND VGND VPWR VPWR _00902_ sky130_fd_sc_hd__mux2_1
XFILLER_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09079_ net970 net3026 net410 VGND VGND VPWR VPWR _00833_ sky130_fd_sc_hd__mux2_1
XFILLER_162_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11110_ net1078 net3801 net543 VGND VGND VPWR VPWR _02853_ sky130_fd_sc_hd__mux2_1
XFILLER_135_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12090_ clknet_leaf_82_clk _00898_ VGND VGND VPWR VPWR data_array.data1\[14\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold770 data_array.data0\[9\]\[5\] VGND VGND VPWR VPWR net2421 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold781 data_array.data1\[5\]\[25\] VGND VGND VPWR VPWR net2432 sky130_fd_sc_hd__dlygate4sd3_1
Xhold792 data_array.data0\[10\]\[2\] VGND VGND VPWR VPWR net2443 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11041_ net2310 net1096 net334 VGND VGND VPWR VPWR _02784_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_183_3867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_183_3878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2160 tag_array.tag1\[14\]\[9\] VGND VGND VPWR VPWR net3811 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2171 data_array.data0\[3\]\[46\] VGND VGND VPWR VPWR net3822 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2182 data_array.data1\[6\]\[52\] VGND VGND VPWR VPWR net3833 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_92_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2193 data_array.data1\[11\]\[1\] VGND VGND VPWR VPWR net3844 sky130_fd_sc_hd__dlygate4sd3_1
X_12992_ clknet_leaf_112_clk _01686_ VGND VGND VPWR VPWR data_array.data0\[3\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1470 data_array.data1\[15\]\[62\] VGND VGND VPWR VPWR net3121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1481 data_array.data1\[13\]\[32\] VGND VGND VPWR VPWR net3132 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1492 tag_array.tag1\[6\]\[22\] VGND VGND VPWR VPWR net3143 sky130_fd_sc_hd__dlygate4sd3_1
X_11943_ clknet_leaf_249_clk _00751_ VGND VGND VPWR VPWR data_array.data0\[4\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_45_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11874_ clknet_leaf_94_clk _00682_ VGND VGND VPWR VPWR data_array.data0\[5\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_13613_ clknet_leaf_88_clk _02242_ VGND VGND VPWR VPWR data_array.data0\[9\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
X_10825_ net1779 net930 net503 VGND VGND VPWR VPWR _02570_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13544_ clknet_leaf_256_clk _02173_ VGND VGND VPWR VPWR data_array.data1\[0\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
X_10756_ net950 net2979 net500 VGND VGND VPWR VPWR _02501_ sky130_fd_sc_hd__mux2_1
XFILLER_9_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13475_ clknet_leaf_180_clk _02105_ VGND VGND VPWR VPWR tag_array.tag0\[15\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_10687_ net3467 net968 net480 VGND VGND VPWR VPWR _02432_ sky130_fd_sc_hd__mux2_1
XFILLER_139_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12426_ clknet_leaf_84_clk _01120_ VGND VGND VPWR VPWR data_array.data0\[14\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_139_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput308 net308 VGND VGND VPWR VPWR mem_wdata[50] sky130_fd_sc_hd__buf_2
Xoutput319 net319 VGND VGND VPWR VPWR mem_wdata[60] sky130_fd_sc_hd__buf_2
XFILLER_153_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12357_ clknet_leaf_253_clk _00032_ VGND VGND VPWR VPWR data_array.rdata0\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_58_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11308_ net1062 net3666 net801 VGND VGND VPWR VPWR _03051_ sky130_fd_sc_hd__mux2_1
X_12288_ clknet_leaf_234_clk _01046_ VGND VGND VPWR VPWR tag_array.tag1\[13\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_142_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14027_ clknet_leaf_28_clk _02656_ VGND VGND VPWR VPWR data_array.data1\[6\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_11239_ net1075 net2474 net681 VGND VGND VPWR VPWR _02982_ sky130_fd_sc_hd__mux2_1
XFILLER_110_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05800_ _03155_ _03157_ VGND VGND VPWR VPWR _03317_ sky130_fd_sc_hd__or2_1
X_06780_ _04080_ _04081_ VGND VGND VPWR VPWR _00033_ sky130_fd_sc_hd__or2_1
XFILLER_49_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_69_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05731_ fsm.tag_out1\[9\] net8 VGND VGND VPWR VPWR _03248_ sky130_fd_sc_hd__and2b_1
XFILLER_82_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_141_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08450_ net2410 net877 net688 VGND VGND VPWR VPWR _00279_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05662_ net15 fsm.tag_out0\[15\] VGND VGND VPWR VPWR _03179_ sky130_fd_sc_hd__and2b_1
XFILLER_36_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07401_ data_array.data0\[13\]\[60\] net1603 net1507 data_array.data0\[14\]\[60\]
+ VGND VGND VPWR VPWR _04646_ sky130_fd_sc_hd__a22o_1
X_08381_ net2226 net971 net686 VGND VGND VPWR VPWR _00256_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_82_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07332_ data_array.data0\[8\]\[54\] net1356 net1262 data_array.data0\[11\]\[54\]
+ _04582_ VGND VGND VPWR VPWR _04583_ sky130_fd_sc_hd__a221o_1
XFILLER_91_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07263_ net1177 _04515_ _04519_ net1225 VGND VGND VPWR VPWR _04521_ sky130_fd_sc_hd__a22o_1
XFILLER_176_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09002_ net2275 net1018 net421 VGND VGND VPWR VPWR _00757_ sky130_fd_sc_hd__mux2_1
X_06214_ tag_array.tag0\[12\]\[2\] net1369 net1275 tag_array.tag0\[15\]\[2\] _03566_
+ VGND VGND VPWR VPWR _03567_ sky130_fd_sc_hd__a221o_1
XFILLER_118_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07194_ data_array.data0\[1\]\[41\] net1529 net1433 data_array.data0\[2\]\[41\] VGND
+ VGND VPWR VPWR _04458_ sky130_fd_sc_hd__a22o_1
X_06145_ data_array.rdata0\[60\] _03477_ _03480_ data_array.rdata1\[60\] VGND VGND
+ VPWR VPWR net319 sky130_fd_sc_hd__a22o_1
XFILLER_145_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_148_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06076_ fsm.tag_out0\[20\] net1120 _03501_ VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__a21o_1
XFILLER_144_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_165_3531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout502 net504 VGND VGND VPWR VPWR net502 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_6_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09904_ net793 net3998 net603 VGND VGND VPWR VPWR _01654_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_6_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout513 _05600_ VGND VGND VPWR VPWR net513 sky130_fd_sc_hd__clkbuf_4
Xfanout524 net525 VGND VGND VPWR VPWR net524 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_165_3542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout535 net537 VGND VGND VPWR VPWR net535 sky130_fd_sc_hd__clkbuf_8
Xfanout546 net547 VGND VGND VPWR VPWR net546 sky130_fd_sc_hd__buf_4
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09835_ net868 net2400 net392 VGND VGND VPWR VPWR _01586_ sky130_fd_sc_hd__mux2_1
Xfanout557 net560 VGND VGND VPWR VPWR net557 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout568 net572 VGND VGND VPWR VPWR net568 sky130_fd_sc_hd__clkbuf_8
XFILLER_112_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout579 net581 VGND VGND VPWR VPWR net579 sky130_fd_sc_hd__clkbuf_4
XFILLER_101_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09766_ net2871 net724 net671 VGND VGND VPWR VPWR _01518_ sky130_fd_sc_hd__mux2_1
XFILLER_6_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06978_ _04260_ _04261_ VGND VGND VPWR VPWR _00013_ sky130_fd_sc_hd__or2_1
XFILLER_39_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08717_ net3680 net756 net475 VGND VGND VPWR VPWR _00476_ sky130_fd_sc_hd__mux2_1
X_05929_ net124 net1150 _03412_ _03413_ VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__a22o_1
XFILLER_73_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09697_ net698 net2834 net606 VGND VGND VPWR VPWR _01449_ sky130_fd_sc_hd__mux2_1
XFILLER_27_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08648_ net2007 net730 net507 VGND VGND VPWR VPWR _00407_ sky130_fd_sc_hd__mux2_1
XFILLER_41_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08579_ net1275 net1199 net814 net1709 VGND VGND VPWR VPWR _00340_ sky130_fd_sc_hd__a31o_1
XFILLER_168_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10610_ net2040 net1022 net467 VGND VGND VPWR VPWR _02355_ sky130_fd_sc_hd__mux2_1
X_11590_ clknet_leaf_195_clk _00398_ VGND VGND VPWR VPWR tag_array.tag1\[4\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_10 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10541_ net1041 net2094 net454 VGND VGND VPWR VPWR _02286_ sky130_fd_sc_hd__mux2_1
XFILLER_155_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13260_ clknet_leaf_89_clk _01890_ VGND VGND VPWR VPWR data_array.data0\[11\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
X_10472_ net1058 net3009 net346 VGND VGND VPWR VPWR _02217_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_137_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Left_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12211_ clknet_leaf_150_clk _00140_ VGND VGND VPWR VPWR fsm.tag_out0\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_109_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13191_ clknet_leaf_14_clk _00084_ VGND VGND VPWR VPWR data_array.rdata1\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_151_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12142_ clknet_leaf_182_clk _00950_ VGND VGND VPWR VPWR tag_array.tag0\[12\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_12073_ clknet_leaf_67_clk _00881_ VGND VGND VPWR VPWR data_array.data1\[14\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11024_ net1805 net904 net336 VGND VGND VPWR VPWR _02768_ sky130_fd_sc_hd__mux2_1
XFILLER_89_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_86_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_32_Left_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12975_ clknet_leaf_165_clk _01669_ VGND VGND VPWR VPWR tag_array.tag0\[4\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_80_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11926_ clknet_leaf_230_clk _00734_ VGND VGND VPWR VPWR data_array.data0\[4\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11857_ clknet_leaf_52_clk _00665_ VGND VGND VPWR VPWR data_array.data0\[7\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
X_10808_ net2028 net997 net504 VGND VGND VPWR VPWR _02553_ sky130_fd_sc_hd__mux2_1
X_11788_ clknet_leaf_222_clk _00596_ VGND VGND VPWR VPWR data_array.data0\[8\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_60_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13527_ clknet_leaf_91_clk _02156_ VGND VGND VPWR VPWR data_array.data1\[0\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_158_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10739_ net1016 net3402 net493 VGND VGND VPWR VPWR _02484_ sky130_fd_sc_hd__mux2_1
XFILLER_9_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_387 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Left_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13458_ clknet_leaf_231_clk _02088_ VGND VGND VPWR VPWR tag_array.tag0\[1\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_174_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12409_ clknet_leaf_237_clk _01103_ VGND VGND VPWR VPWR data_array.data0\[14\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_127_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13389_ clknet_leaf_57_clk _02019_ VGND VGND VPWR VPWR data_array.data1\[8\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_58_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07950_ data_array.data1\[4\]\[46\] net1333 net1239 data_array.data1\[7\]\[46\] _05144_
+ VGND VGND VPWR VPWR _05145_ sky130_fd_sc_hd__a221o_1
Xhold2907 data_array.data0\[11\]\[3\] VGND VGND VPWR VPWR net4558 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_141_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2918 data_array.data1\[10\]\[28\] VGND VGND VPWR VPWR net4569 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2929 data_array.data0\[15\]\[30\] VGND VGND VPWR VPWR net4580 sky130_fd_sc_hd__dlygate4sd3_1
X_06901_ _04190_ _04191_ VGND VGND VPWR VPWR _00005_ sky130_fd_sc_hd__or2_1
X_07881_ data_array.data1\[13\]\[40\] net1606 net1510 data_array.data1\[14\]\[40\]
+ VGND VGND VPWR VPWR _05082_ sky130_fd_sc_hd__a22o_1
XFILLER_122_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_143_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09620_ net868 net4249 net400 VGND VGND VPWR VPWR _01372_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_50_Left_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06832_ data_array.data0\[0\]\[8\] net1345 net1251 data_array.data0\[3\]\[8\] _04128_
+ VGND VGND VPWR VPWR _04129_ sky130_fd_sc_hd__a221o_1
XFILLER_37_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09551_ net723 net3706 net619 VGND VGND VPWR VPWR _01304_ sky130_fd_sc_hd__mux2_1
XFILLER_37_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06763_ data_array.data0\[9\]\[2\] net1528 net1432 data_array.data0\[10\]\[2\] VGND
+ VGND VPWR VPWR _04066_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_121_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08502_ net1720 net617 VGND VGND VPWR VPWR _00296_ sky130_fd_sc_hd__nand2b_1
XFILLER_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05714_ _03227_ _03228_ _03230_ VGND VGND VPWR VPWR _03231_ sky130_fd_sc_hd__or3_1
X_09482_ net700 net4158 net659 VGND VGND VPWR VPWR _01235_ sky130_fd_sc_hd__mux2_1
XFILLER_52_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06694_ tag_array.tag1\[8\]\[21\] net1401 net1307 tag_array.tag1\[11\]\[21\] _04002_
+ VGND VGND VPWR VPWR _04003_ sky130_fd_sc_hd__a221o_1
X_08433_ net147 net82 net1638 VGND VGND VPWR VPWR _05525_ sky130_fd_sc_hd__mux2_1
X_05645_ _03160_ _03161_ fsm.valid0 VGND VGND VPWR VPWR _03162_ sky130_fd_sc_hd__or3b_1
XFILLER_24_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08364_ net122 net57 net1641 VGND VGND VPWR VPWR _05479_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07315_ data_array.data0\[1\]\[52\] net1548 net1452 data_array.data0\[2\]\[52\] VGND
+ VGND VPWR VPWR _04568_ sky130_fd_sc_hd__a22o_1
X_08295_ net160 net95 net1641 VGND VGND VPWR VPWR _05433_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_119_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07246_ data_array.data0\[4\]\[46\] net1341 net1247 data_array.data0\[7\]\[46\] _04504_
+ VGND VGND VPWR VPWR _04505_ sky130_fd_sc_hd__a221o_1
XFILLER_176_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_335 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07177_ data_array.data0\[13\]\[40\] net1602 net1506 data_array.data0\[14\]\[40\]
+ VGND VGND VPWR VPWR _04442_ sky130_fd_sc_hd__a22o_1
XFILLER_11_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06128_ data_array.rdata0\[43\] net1140 net1114 data_array.rdata1\[43\] VGND VGND
+ VPWR VPWR net300 sky130_fd_sc_hd__a22o_1
X_06059_ net1159 net11 fsm.tag_out1\[12\] net1131 VGND VGND VPWR VPWR _03493_ sky130_fd_sc_hd__a22o_1
Xfanout1308 net1309 VGND VGND VPWR VPWR net1308 sky130_fd_sc_hd__clkbuf_4
Xfanout1319 net1328 VGND VGND VPWR VPWR net1319 sky130_fd_sc_hd__clkbuf_4
Xfanout332 _03133_ VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_180_3815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout343 _03132_ VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__buf_4
XFILLER_115_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_180_3826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout354 net355 VGND VGND VPWR VPWR net354 sky130_fd_sc_hd__buf_4
Xfanout365 net369 VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__clkbuf_4
Xfanout376 _03127_ VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__buf_4
Xfanout387 net393 VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__clkbuf_8
X_09818_ net939 net3498 net390 VGND VGND VPWR VPWR _01569_ sky130_fd_sc_hd__mux2_1
XFILLER_115_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout398 net400 VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__clkbuf_8
XFILLER_98_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09749_ net1807 net791 net667 VGND VGND VPWR VPWR _01501_ sky130_fd_sc_hd__mux2_1
X_12760_ clknet_leaf_177_clk _01454_ VGND VGND VPWR VPWR tag_array.tag0\[6\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_178_3777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11711_ clknet_leaf_170_clk _00519_ VGND VGND VPWR VPWR tag_array.tag0\[9\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_178_3788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ clknet_leaf_158_clk _01385_ VGND VGND VPWR VPWR tag_array.tag0\[8\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_159_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14430_ clknet_leaf_42_clk _03053_ VGND VGND VPWR VPWR data_array.data1\[7\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_42_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11642_ clknet_leaf_139_clk _00450_ VGND VGND VPWR VPWR tag_array.tag1\[2\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_14361_ clknet_leaf_34_clk _02984_ VGND VGND VPWR VPWR data_array.data1\[10\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11573_ clknet_leaf_232_clk _00381_ VGND VGND VPWR VPWR tag_array.tag1\[5\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput18 cpu_addr[25] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_2
X_13312_ clknet_leaf_228_clk _01942_ VGND VGND VPWR VPWR data_array.data0\[10\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10524_ net1111 net2798 net458 VGND VGND VPWR VPWR _02269_ sky130_fd_sc_hd__mux2_1
Xinput29 cpu_addr[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_4
XFILLER_182_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14292_ clknet_leaf_84_clk _02921_ VGND VGND VPWR VPWR data_array.data1\[11\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_155_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13243_ clknet_leaf_224_clk _01873_ VGND VGND VPWR VPWR data_array.data0\[11\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_182_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10455_ net2568 net352 net479 VGND VGND VPWR VPWR _02201_ sky130_fd_sc_hd__mux2_1
XFILLER_6_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13174_ clknet_leaf_49_clk _00066_ VGND VGND VPWR VPWR data_array.rdata1\[11\] sky130_fd_sc_hd__dfxtp_1
X_10386_ net2096 net1110 net665 VGND VGND VPWR VPWR _02132_ sky130_fd_sc_hd__mux2_1
XFILLER_124_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_107_Left_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12125_ clknet_leaf_144_clk _00933_ VGND VGND VPWR VPWR tag_array.tag0\[12\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_176_Right_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12056_ clknet_leaf_251_clk _00864_ VGND VGND VPWR VPWR data_array.data1\[14\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_111_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11007_ net2128 net972 net336 VGND VGND VPWR VPWR _02751_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12958_ clknet_leaf_110_clk _01652_ VGND VGND VPWR VPWR data_array.data0\[13\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
X_11909_ clknet_leaf_90_clk _00717_ VGND VGND VPWR VPWR data_array.data0\[5\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
X_12889_ clknet_leaf_234_clk _01583_ VGND VGND VPWR VPWR data_array.data0\[12\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_16_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07100_ data_array.data0\[13\]\[33\] net1585 net1489 data_array.data0\[14\]\[33\]
+ VGND VGND VPWR VPWR _04372_ sky130_fd_sc_hd__a22o_1
X_08080_ data_array.data1\[8\]\[58\] net1359 net1265 data_array.data1\[11\]\[58\]
+ _05262_ VGND VGND VPWR VPWR _05263_ sky130_fd_sc_hd__a221o_1
Xclkload201 clknet_leaf_164_clk VGND VGND VPWR VPWR clkload201/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload212 clknet_leaf_120_clk VGND VGND VPWR VPWR clkload212/X sky130_fd_sc_hd__clkbuf_8
X_07031_ net1617 _04303_ _04307_ net1191 VGND VGND VPWR VPWR _04310_ sky130_fd_sc_hd__a22o_1
Xclkload223 clknet_leaf_162_clk VGND VGND VPWR VPWR clkload223/Y sky130_fd_sc_hd__bufinv_16
Xclkload234 clknet_leaf_132_clk VGND VGND VPWR VPWR clkload234/Y sky130_fd_sc_hd__inv_8
XFILLER_134_508 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload245 clknet_leaf_146_clk VGND VGND VPWR VPWR clkload245/Y sky130_fd_sc_hd__inv_8
XFILLER_174_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_263_clk clknet_5_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_263_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_142_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08982_ net2178 net1096 net423 VGND VGND VPWR VPWR _00737_ sky130_fd_sc_hd__mux2_1
Xhold2704 tag_array.tag1\[5\]\[1\] VGND VGND VPWR VPWR net4355 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_143_Right_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2715 data_array.data1\[9\]\[51\] VGND VGND VPWR VPWR net4366 sky130_fd_sc_hd__dlygate4sd3_1
X_07933_ net1631 _05123_ _05127_ net1205 VGND VGND VPWR VPWR _05130_ sky130_fd_sc_hd__a22o_1
Xhold2726 data_array.data0\[13\]\[41\] VGND VGND VPWR VPWR net4377 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_110_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2737 data_array.data0\[13\]\[47\] VGND VGND VPWR VPWR net4388 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2748 tag_array.tag0\[15\]\[15\] VGND VGND VPWR VPWR net4399 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2759 data_array.data1\[6\]\[1\] VGND VGND VPWR VPWR net4410 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07864_ data_array.data1\[12\]\[38\] net1398 net1304 data_array.data1\[15\]\[38\]
+ _05066_ VGND VGND VPWR VPWR _05067_ sky130_fd_sc_hd__a221o_1
XFILLER_69_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09603_ net936 net3600 net398 VGND VGND VPWR VPWR _01355_ sky130_fd_sc_hd__mux2_1
XFILLER_113_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06815_ data_array.data0\[8\]\[7\] net1395 net1301 data_array.data0\[11\]\[7\] _04112_
+ VGND VGND VPWR VPWR _04113_ sky130_fd_sc_hd__a221o_1
X_07795_ data_array.data1\[1\]\[32\] net1520 net1424 data_array.data1\[2\]\[32\] VGND
+ VGND VPWR VPWR _05004_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_27_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09534_ net793 net2732 net619 VGND VGND VPWR VPWR _01287_ sky130_fd_sc_hd__mux2_1
X_06746_ net1222 _04045_ _04049_ net1173 VGND VGND VPWR VPWR _04051_ sky130_fd_sc_hd__a22o_1
XFILLER_71_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09465_ net767 net4117 net653 VGND VGND VPWR VPWR _01218_ sky130_fd_sc_hd__mux2_1
X_06677_ tag_array.tag1\[1\]\[19\] net1592 net1496 tag_array.tag1\[2\]\[19\] VGND
+ VGND VPWR VPWR _03988_ sky130_fd_sc_hd__a22o_1
XFILLER_19_1028 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08416_ net1128 _05513_ VGND VGND VPWR VPWR _05514_ sky130_fd_sc_hd__and2_2
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05628_ net1644 net33 VGND VGND VPWR VPWR _03148_ sky130_fd_sc_hd__nor2_1
X_09396_ net1082 net2691 net587 VGND VGND VPWR VPWR _01149_ sky130_fd_sc_hd__mux2_1
XFILLER_145_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08347_ net1127 _05467_ VGND VGND VPWR VPWR _05468_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_173_3685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08278_ net1124 _05421_ VGND VGND VPWR VPWR _05422_ sky130_fd_sc_hd__and2_1
XFILLER_138_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07229_ net1632 _04483_ _04487_ net1206 VGND VGND VPWR VPWR _04490_ sky130_fd_sc_hd__a22o_1
XFILLER_164_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10240_ net784 net4053 net595 VGND VGND VPWR VPWR _01987_ sky130_fd_sc_hd__mux2_1
XFILLER_3_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_254_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_254_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10171_ net861 net2337 net369 VGND VGND VPWR VPWR _01919_ sky130_fd_sc_hd__mux2_1
Xfanout1105 net1106 VGND VGND VPWR VPWR net1105 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_110_Right_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1116 _03480_ VGND VGND VPWR VPWR net1116 sky130_fd_sc_hd__buf_8
XFILLER_120_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1127 net1128 VGND VGND VPWR VPWR net1127 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1138 _03477_ VGND VGND VPWR VPWR net1138 sky130_fd_sc_hd__clkbuf_8
Xfanout1149 _03154_ VGND VGND VPWR VPWR net1149 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_35_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13930_ clknet_leaf_8_clk _02559_ VGND VGND VPWR VPWR data_array.data1\[4\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13861_ clknet_leaf_40_clk _02490_ VGND VGND VPWR VPWR data_array.data1\[3\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_170_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12812_ clknet_leaf_135_clk _01506_ VGND VGND VPWR VPWR tag_array.tag1\[0\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_13792_ clknet_leaf_91_clk _02421_ VGND VGND VPWR VPWR data_array.data1\[2\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12743_ clknet_leaf_166_clk _01437_ VGND VGND VPWR VPWR tag_array.tag0\[5\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12674_ clknet_leaf_13_clk _01368_ VGND VGND VPWR VPWR data_array.data0\[15\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
X_14413_ clknet_leaf_192_clk _03036_ VGND VGND VPWR VPWR data_array.data1\[10\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
X_11625_ clknet_leaf_140_clk _00433_ VGND VGND VPWR VPWR tag_array.tag1\[3\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_13_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14344_ clknet_leaf_184_clk _00186_ _00189_ VGND VGND VPWR VPWR fsm.state\[0\] sky130_fd_sc_hd__dfstp_1
XFILLER_184_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11556_ clknet_leaf_194_clk _00364_ VGND VGND VPWR VPWR tag_array.tag1\[6\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_156_666 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10507_ net917 net3354 net349 VGND VGND VPWR VPWR _02252_ sky130_fd_sc_hd__mux2_1
X_14275_ clknet_leaf_41_clk _02904_ VGND VGND VPWR VPWR data_array.data1\[12\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_156_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11487_ clknet_leaf_151_clk _00296_ VGND VGND VPWR VPWR tag_array.valid0\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_137_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_115_Left_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13226_ clknet_leaf_202_clk _00123_ VGND VGND VPWR VPWR data_array.rdata1\[63\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_94_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10438_ net2484 net900 net664 VGND VGND VPWR VPWR _02184_ sky130_fd_sc_hd__mux2_1
XFILLER_170_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_245_clk clknet_5_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_245_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_55_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13157_ clknet_leaf_103_clk _01851_ VGND VGND VPWR VPWR tag_array.tag1\[8\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_10369_ net723 net2939 net539 VGND VGND VPWR VPWR _02116_ sky130_fd_sc_hd__mux2_1
X_12108_ clknet_leaf_251_clk _00916_ VGND VGND VPWR VPWR data_array.data1\[14\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_72_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13088_ clknet_leaf_240_clk _01782_ VGND VGND VPWR VPWR data_array.data1\[13\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_72_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1650 net1651 VGND VGND VPWR VPWR net1650 sky130_fd_sc_hd__clkbuf_2
X_12039_ clknet_leaf_53_clk _00847_ VGND VGND VPWR VPWR data_array.data0\[6\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_1_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_1_0_clk sky130_fd_sc_hd__clkbuf_8
X_06600_ tag_array.tag1\[1\]\[12\] net1592 net1496 tag_array.tag1\[2\]\[12\] VGND
+ VGND VPWR VPWR _03918_ sky130_fd_sc_hd__a22o_1
XFILLER_19_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07580_ data_array.data1\[4\]\[12\] net1395 net1301 data_array.data1\[7\]\[12\] _04808_
+ VGND VGND VPWR VPWR _04809_ sky130_fd_sc_hd__a221o_1
X_06531_ tag_array.tag1\[0\]\[6\] net1362 net1268 tag_array.tag1\[3\]\[6\] _03854_
+ VGND VGND VPWR VPWR _03855_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_138_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09250_ net779 net4566 net571 VGND VGND VPWR VPWR _01004_ sky130_fd_sc_hd__mux2_1
X_06462_ tag_array.tag1\[9\]\[0\] net1591 net1495 tag_array.tag1\[10\]\[0\] VGND VGND
+ VPWR VPWR _03792_ sky130_fd_sc_hd__a22o_1
XFILLER_167_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08201_ fsm.tag_out1\[2\] net816 net808 fsm.tag_out0\[2\] _05368_ VGND VGND VPWR
+ VPWR _05369_ sky130_fd_sc_hd__a221o_4
XFILLER_18_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06393_ net1201 _03723_ _03727_ net1626 VGND VGND VPWR VPWR _03730_ sky130_fd_sc_hd__a22o_1
X_09181_ net755 net2539 net628 VGND VGND VPWR VPWR _00935_ sky130_fd_sc_hd__mux2_1
XFILLER_159_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08132_ net1183 _05305_ _05309_ net1233 VGND VGND VPWR VPWR _05311_ sky130_fd_sc_hd__a22o_1
XFILLER_175_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08063_ data_array.data1\[1\]\[56\] net1533 net1437 data_array.data1\[2\]\[56\] VGND
+ VGND VPWR VPWR _05248_ sky130_fd_sc_hd__a22o_1
XFILLER_88_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07014_ data_array.data0\[1\]\[25\] net1519 net1423 data_array.data0\[2\]\[25\] VGND
+ VGND VPWR VPWR _04294_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_112_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_236_clk clknet_5_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_236_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_382 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_747 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2501 tag_array.tag0\[15\]\[13\] VGND VGND VPWR VPWR net4152 sky130_fd_sc_hd__dlygate4sd3_1
X_08965_ net904 net3230 net426 VGND VGND VPWR VPWR _00721_ sky130_fd_sc_hd__mux2_1
Xhold2512 tag_array.tag1\[3\]\[3\] VGND VGND VPWR VPWR net4163 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2523 data_array.data1\[6\]\[38\] VGND VGND VPWR VPWR net4174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2534 data_array.data1\[15\]\[4\] VGND VGND VPWR VPWR net4185 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1800 tag_array.tag1\[14\]\[5\] VGND VGND VPWR VPWR net3451 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2545 data_array.data0\[14\]\[21\] VGND VGND VPWR VPWR net4196 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2556 data_array.data1\[11\]\[30\] VGND VGND VPWR VPWR net4207 sky130_fd_sc_hd__dlygate4sd3_1
X_07916_ data_array.data1\[1\]\[43\] net1568 net1472 data_array.data1\[2\]\[43\] VGND
+ VGND VPWR VPWR _05114_ sky130_fd_sc_hd__a22o_1
Xhold1811 tag_array.tag0\[4\]\[10\] VGND VGND VPWR VPWR net3462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1822 data_array.data1\[9\]\[56\] VGND VGND VPWR VPWR net3473 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_25_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2567 data_array.data1\[6\]\[51\] VGND VGND VPWR VPWR net4218 sky130_fd_sc_hd__dlygate4sd3_1
X_08896_ net921 net3640 net439 VGND VGND VPWR VPWR _00653_ sky130_fd_sc_hd__mux2_1
Xhold1833 tag_array.tag1\[3\]\[22\] VGND VGND VPWR VPWR net3484 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2578 data_array.data0\[3\]\[49\] VGND VGND VPWR VPWR net4229 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2589 data_array.data1\[6\]\[25\] VGND VGND VPWR VPWR net4240 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1844 data_array.data1\[12\]\[39\] VGND VGND VPWR VPWR net3495 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1855 data_array.data1\[14\]\[12\] VGND VGND VPWR VPWR net3506 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07847_ _05050_ _05051_ VGND VGND VPWR VPWR _00093_ sky130_fd_sc_hd__or2_1
Xhold1866 data_array.data0\[12\]\[46\] VGND VGND VPWR VPWR net3517 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1877 data_array.data0\[11\]\[61\] VGND VGND VPWR VPWR net3528 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1888 data_array.data0\[13\]\[13\] VGND VGND VPWR VPWR net3539 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1899 data_array.data0\[15\]\[52\] VGND VGND VPWR VPWR net3550 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_95_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07778_ data_array.data1\[0\]\[30\] net1400 net1306 data_array.data1\[3\]\[30\] _04988_
+ VGND VGND VPWR VPWR _04989_ sky130_fd_sc_hd__a221o_1
X_09517_ net761 net3395 net623 VGND VGND VPWR VPWR _01270_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_175_3714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06729_ tag_array.tag1\[4\]\[24\] net1372 net1278 tag_array.tag1\[7\]\[24\] _04034_
+ VGND VGND VPWR VPWR _04035_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_175_3725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09448_ net874 net2852 net585 VGND VGND VPWR VPWR _01201_ sky130_fd_sc_hd__mux2_1
XFILLER_13_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09379_ net885 net2366 net403 VGND VGND VPWR VPWR _01132_ sky130_fd_sc_hd__mux2_1
XFILLER_8_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11410_ clknet_leaf_189_clk _00220_ VGND VGND VPWR VPWR tag_array.tag1\[7\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_137_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12390_ clknet_leaf_16_clk _01084_ VGND VGND VPWR VPWR data_array.data0\[14\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11341_ net930 net3415 net796 VGND VGND VPWR VPWR _03084_ sky130_fd_sc_hd__mux2_1
XFILLER_126_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14060_ clknet_leaf_82_clk _02689_ VGND VGND VPWR VPWR data_array.data1\[6\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
X_11272_ net943 net4137 net682 VGND VGND VPWR VPWR _03015_ sky130_fd_sc_hd__mux2_1
XFILLER_4_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13011_ clknet_leaf_246_clk _01705_ VGND VGND VPWR VPWR data_array.data0\[3\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_227_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_227_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10223_ net913 net2050 net359 VGND VGND VPWR VPWR _01970_ sky130_fd_sc_hd__mux2_1
XFILLER_121_522 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10154_ net929 net3868 net363 VGND VGND VPWR VPWR _01902_ sky130_fd_sc_hd__mux2_1
XFILLER_66_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10085_ net1822 net783 net636 VGND VGND VPWR VPWR _01834_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13913_ clknet_leaf_253_clk _02542_ VGND VGND VPWR VPWR data_array.data1\[4\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13844_ clknet_leaf_85_clk _02473_ VGND VGND VPWR VPWR data_array.data1\[3\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_18_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13775_ clknet_leaf_83_clk _02404_ VGND VGND VPWR VPWR data_array.data1\[2\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_10987_ net2603 net1052 net342 VGND VGND VPWR VPWR _02731_ sky130_fd_sc_hd__mux2_1
XFILLER_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12726_ clknet_leaf_106_clk _01420_ VGND VGND VPWR VPWR tag_array.tag0\[7\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_745 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12657_ clknet_leaf_234_clk _01351_ VGND VGND VPWR VPWR data_array.data0\[15\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_88_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_96_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11608_ clknet_leaf_188_clk _00416_ VGND VGND VPWR VPWR tag_array.tag1\[4\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_96_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12588_ clknet_leaf_169_clk _01282_ VGND VGND VPWR VPWR tag_array.tag0\[10\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_157_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14327_ clknet_leaf_79_clk _02956_ VGND VGND VPWR VPWR data_array.data1\[11\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
X_11539_ clknet_leaf_129_clk _00347_ VGND VGND VPWR VPWR tag_array.tag1\[6\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold407 data_array.data1\[2\]\[34\] VGND VGND VPWR VPWR net2058 sky130_fd_sc_hd__dlygate4sd3_1
Xhold418 tag_array.tag0\[8\]\[21\] VGND VGND VPWR VPWR net2069 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14258_ clknet_leaf_84_clk _02887_ VGND VGND VPWR VPWR data_array.data1\[12\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold429 tag_array.tag0\[3\]\[21\] VGND VGND VPWR VPWR net2080 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_218_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_218_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_98_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13209_ clknet_leaf_266_clk _00104_ VGND VGND VPWR VPWR data_array.rdata1\[46\] sky130_fd_sc_hd__dfxtp_1
X_14189_ clknet_leaf_218_clk _02818_ VGND VGND VPWR VPWR data_array.data0\[2\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout909 net910 VGND VGND VPWR VPWR net909 sky130_fd_sc_hd__clkbuf_2
XFILLER_97_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08750_ net725 net3412 net463 VGND VGND VPWR VPWR _00509_ sky130_fd_sc_hd__mux2_1
Xhold1107 tag_array.tag0\[10\]\[5\] VGND VGND VPWR VPWR net2758 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1118 data_array.data0\[5\]\[39\] VGND VGND VPWR VPWR net2769 sky130_fd_sc_hd__dlygate4sd3_1
X_05962_ net136 net1156 _03434_ _03435_ VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__a22o_1
Xhold1129 data_array.data0\[6\]\[52\] VGND VGND VPWR VPWR net2780 sky130_fd_sc_hd__dlygate4sd3_1
X_07701_ data_array.data1\[4\]\[23\] net1360 net1266 data_array.data1\[7\]\[23\] _04918_
+ VGND VGND VPWR VPWR _04919_ sky130_fd_sc_hd__a221o_1
Xfanout1480 net1495 VGND VGND VPWR VPWR net1480 sky130_fd_sc_hd__clkbuf_4
X_08681_ net701 net3112 net501 VGND VGND VPWR VPWR _00440_ sky130_fd_sc_hd__mux2_1
Xfanout1491 net1495 VGND VGND VPWR VPWR net1491 sky130_fd_sc_hd__clkbuf_2
X_05893_ net111 net1157 _03388_ _03389_ VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__a22o_1
X_07632_ data_array.data1\[9\]\[17\] net1526 net1430 data_array.data1\[10\]\[17\]
+ VGND VGND VPWR VPWR _04856_ sky130_fd_sc_hd__a22o_1
XFILLER_54_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07563_ data_array.data1\[8\]\[11\] net1385 net1291 data_array.data1\[11\]\[11\]
+ _04792_ VGND VGND VPWR VPWR _04793_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_105_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09302_ net772 net2524 net551 VGND VGND VPWR VPWR _01056_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06514_ net1623 _03833_ _03837_ net1197 VGND VGND VPWR VPWR _03840_ sky130_fd_sc_hd__a22o_1
XFILLER_181_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07494_ net1178 _04725_ _04729_ net1226 VGND VGND VPWR VPWR _04731_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_153_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09233_ net749 net3904 net645 VGND VGND VPWR VPWR _00987_ sky130_fd_sc_hd__mux2_1
XFILLER_181_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_588 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06445_ tag_array.tag0\[12\]\[23\] net1409 net1315 tag_array.tag0\[15\]\[23\] _03776_
+ VGND VGND VPWR VPWR _03777_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_170_3622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09164_ net886 net4395 net568 VGND VGND VPWR VPWR _00918_ sky130_fd_sc_hd__mux2_1
X_06376_ tag_array.tag0\[5\]\[17\] net1602 net1506 tag_array.tag0\[6\]\[17\] VGND
+ VGND VPWR VPWR _03714_ sky130_fd_sc_hd__a22o_1
XFILLER_163_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08115_ data_array.data1\[0\]\[61\] net1359 net1265 data_array.data1\[3\]\[61\] _05294_
+ VGND VGND VPWR VPWR _05295_ sky130_fd_sc_hd__a221o_1
XFILLER_181_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09095_ net904 net4138 net410 VGND VGND VPWR VPWR _00849_ sky130_fd_sc_hd__mux2_1
X_08046_ data_array.data1\[13\]\[55\] net1535 net1439 data_array.data1\[14\]\[55\]
+ VGND VGND VPWR VPWR _05232_ sky130_fd_sc_hd__a22o_1
XFILLER_31_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold930 data_array.data1\[1\]\[0\] VGND VGND VPWR VPWR net2581 sky130_fd_sc_hd__dlygate4sd3_1
Xhold941 tag_array.tag0\[14\]\[4\] VGND VGND VPWR VPWR net2592 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_209_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_209_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold952 data_array.data0\[1\]\[14\] VGND VGND VPWR VPWR net2603 sky130_fd_sc_hd__dlygate4sd3_1
Xhold963 tag_array.tag0\[12\]\[16\] VGND VGND VPWR VPWR net2614 sky130_fd_sc_hd__dlygate4sd3_1
Xhold974 data_array.data1\[1\]\[28\] VGND VGND VPWR VPWR net2625 sky130_fd_sc_hd__dlygate4sd3_1
Xhold985 tag_array.tag1\[14\]\[6\] VGND VGND VPWR VPWR net2636 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_3584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold996 data_array.data0\[15\]\[61\] VGND VGND VPWR VPWR net2647 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_168_3595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09997_ net1099 net3133 net556 VGND VGND VPWR VPWR _01746_ sky130_fd_sc_hd__mux2_1
Xhold2320 data_array.data1\[15\]\[27\] VGND VGND VPWR VPWR net3971 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2331 data_array.data0\[10\]\[47\] VGND VGND VPWR VPWR net3982 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2342 data_array.data1\[13\]\[40\] VGND VGND VPWR VPWR net3993 sky130_fd_sc_hd__dlygate4sd3_1
X_08948_ net972 net2651 net427 VGND VGND VPWR VPWR _00704_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2353 data_array.data1\[7\]\[18\] VGND VGND VPWR VPWR net4004 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2364 data_array.data1\[7\]\[32\] VGND VGND VPWR VPWR net4015 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1630 data_array.data0\[10\]\[54\] VGND VGND VPWR VPWR net3281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2375 data_array.data1\[15\]\[32\] VGND VGND VPWR VPWR net4026 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1641 data_array.data1\[11\]\[11\] VGND VGND VPWR VPWR net3292 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2386 tag_array.tag1\[13\]\[8\] VGND VGND VPWR VPWR net4037 sky130_fd_sc_hd__dlygate4sd3_1
X_08879_ net988 net4178 net438 VGND VGND VPWR VPWR _00636_ sky130_fd_sc_hd__mux2_1
Xhold2397 tag_array.tag1\[10\]\[8\] VGND VGND VPWR VPWR net4048 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1652 data_array.data0\[14\]\[25\] VGND VGND VPWR VPWR net3303 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1663 data_array.data1\[3\]\[39\] VGND VGND VPWR VPWR net3314 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1674 data_array.data0\[8\]\[13\] VGND VGND VPWR VPWR net3325 sky130_fd_sc_hd__dlygate4sd3_1
X_10910_ net1100 net3590 net527 VGND VGND VPWR VPWR _02655_ sky130_fd_sc_hd__mux2_1
XFILLER_44_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1685 tag_array.tag0\[2\]\[11\] VGND VGND VPWR VPWR net3336 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1696 data_array.data0\[13\]\[4\] VGND VGND VPWR VPWR net3347 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11890_ clknet_leaf_25_clk _00698_ VGND VGND VPWR VPWR data_array.data0\[5\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_10841_ net3070 net864 net506 VGND VGND VPWR VPWR _02586_ sky130_fd_sc_hd__mux2_1
X_13560_ clknet_leaf_248_clk _02189_ VGND VGND VPWR VPWR data_array.data1\[0\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
X_10772_ net886 net3595 net492 VGND VGND VPWR VPWR _02517_ sky130_fd_sc_hd__mux2_1
XFILLER_40_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12511_ clknet_leaf_192_clk _01205_ VGND VGND VPWR VPWR data_array.data1\[9\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
X_13491_ clknet_leaf_182_clk _02121_ VGND VGND VPWR VPWR tag_array.tag0\[15\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_40_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12442_ clknet_leaf_114_clk _01136_ VGND VGND VPWR VPWR data_array.data0\[14\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_139_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12373_ clknet_leaf_14_clk _00050_ VGND VGND VPWR VPWR data_array.rdata0\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14112_ clknet_leaf_92_clk _02741_ VGND VGND VPWR VPWR data_array.data0\[1\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11324_ net997 net4490 net796 VGND VGND VPWR VPWR _03067_ sky130_fd_sc_hd__mux2_1
XFILLER_176_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_1019 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14043_ clknet_leaf_66_clk _02672_ VGND VGND VPWR VPWR data_array.data1\[6\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_141_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11255_ net1008 net3094 net673 VGND VGND VPWR VPWR _02998_ sky130_fd_sc_hd__mux2_1
XFILLER_107_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10206_ net982 net4193 net354 VGND VGND VPWR VPWR _01953_ sky130_fd_sc_hd__mux2_1
XFILLER_79_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11186_ net1031 net3565 net658 VGND VGND VPWR VPWR _02929_ sky130_fd_sc_hd__mux2_1
XFILLER_0_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10137_ net998 net4400 net363 VGND VGND VPWR VPWR _01885_ sky130_fd_sc_hd__mux2_1
XFILLER_94_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10068_ net751 net2582 net600 VGND VGND VPWR VPWR _01817_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_89_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13827_ clknet_leaf_55_clk _02456_ VGND VGND VPWR VPWR data_array.data1\[2\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13758_ clknet_leaf_215_clk _02387_ VGND VGND VPWR VPWR data_array.data1\[1\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12709_ clknet_leaf_168_clk _01403_ VGND VGND VPWR VPWR tag_array.tag0\[7\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_176_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13689_ clknet_leaf_56_clk _02318_ VGND VGND VPWR VPWR data_array.data1\[15\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06230_ _03580_ _03581_ VGND VGND VPWR VPWR _00149_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1042 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06161_ net28 net29 VGND VGND VPWR VPWR _03518_ sky130_fd_sc_hd__nor2_1
XFILLER_184_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_720 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold204 tag_array.tag1\[8\]\[13\] VGND VGND VPWR VPWR net1855 sky130_fd_sc_hd__dlygate4sd3_1
X_06092_ data_array.rdata0\[7\] net1140 net1116 data_array.rdata1\[7\] VGND VGND VPWR
+ VPWR net324 sky130_fd_sc_hd__a22o_1
Xhold215 data_array.data0\[0\]\[59\] VGND VGND VPWR VPWR net1866 sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 data_array.data0\[4\]\[5\] VGND VGND VPWR VPWR net1877 sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 tag_array.tag1\[1\]\[0\] VGND VGND VPWR VPWR net1888 sky130_fd_sc_hd__dlygate4sd3_1
Xhold248 data_array.data0\[8\]\[37\] VGND VGND VPWR VPWR net1899 sky130_fd_sc_hd__dlygate4sd3_1
X_09920_ net727 net3340 net604 VGND VGND VPWR VPWR _01670_ sky130_fd_sc_hd__mux2_1
XFILLER_144_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold259 data_array.data0\[1\]\[24\] VGND VGND VPWR VPWR net1910 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_125_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout706 net707 VGND VGND VPWR VPWR net706 sky130_fd_sc_hd__clkbuf_2
X_09851_ net1064 net2851 net382 VGND VGND VPWR VPWR _01601_ sky130_fd_sc_hd__mux2_1
Xfanout717 _05403_ VGND VGND VPWR VPWR net717 sky130_fd_sc_hd__buf_2
Xfanout728 net729 VGND VGND VPWR VPWR net728 sky130_fd_sc_hd__clkbuf_2
Xfanout739 _05391_ VGND VGND VPWR VPWR net739 sky130_fd_sc_hd__buf_1
XFILLER_140_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08802_ net2173 net1038 net443 VGND VGND VPWR VPWR _00560_ sky130_fd_sc_hd__mux2_1
XFILLER_98_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_146_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09782_ net1080 net2197 net392 VGND VGND VPWR VPWR _01533_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_146_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06994_ data_array.data0\[9\]\[23\] net1561 net1465 data_array.data0\[10\]\[23\]
+ VGND VGND VPWR VPWR _04276_ sky130_fd_sc_hd__a22o_1
XFILLER_22_1013 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08733_ net792 net4108 net460 VGND VGND VPWR VPWR _00492_ sky130_fd_sc_hd__mux2_1
X_05945_ data_array.rdata0\[38\] net1666 net1147 VGND VGND VPWR VPWR _03424_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_163_3492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_1_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08664_ net766 net2793 net493 VGND VGND VPWR VPWR _00423_ sky130_fd_sc_hd__mux2_1
X_05876_ data_array.rdata0\[15\] net850 net1147 VGND VGND VPWR VPWR _03378_ sky130_fd_sc_hd__o21a_1
XFILLER_26_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_124_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07615_ net1180 _04835_ _04839_ net1228 VGND VGND VPWR VPWR _04841_ sky130_fd_sc_hd__a22o_1
X_08595_ net743 net3425 net537 VGND VGND VPWR VPWR _00354_ sky130_fd_sc_hd__mux2_1
XFILLER_179_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07546_ data_array.data1\[1\]\[9\] net1580 net1484 data_array.data1\[2\]\[9\] VGND
+ VGND VPWR VPWR _04778_ sky130_fd_sc_hd__a22o_1
XFILLER_167_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07477_ data_array.data1\[4\]\[3\] net1350 net1256 data_array.data1\[7\]\[3\] _04714_
+ VGND VGND VPWR VPWR _04715_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09216_ net717 net4554 net631 VGND VGND VPWR VPWR _00970_ sky130_fd_sc_hd__mux2_1
X_06428_ _03760_ _03761_ VGND VGND VPWR VPWR _00144_ sky130_fd_sc_hd__or2_1
XFILLER_167_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09147_ net953 net3999 net569 VGND VGND VPWR VPWR _00901_ sky130_fd_sc_hd__mux2_1
X_06359_ tag_array.tag0\[4\]\[15\] net1403 net1309 tag_array.tag0\[7\]\[15\] _03698_
+ VGND VGND VPWR VPWR _03699_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_20_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09078_ net972 net3812 net411 VGND VGND VPWR VPWR _00832_ sky130_fd_sc_hd__mux2_1
XFILLER_136_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08029_ data_array.data1\[12\]\[53\] net1334 net1240 data_array.data1\[15\]\[53\]
+ _05216_ VGND VGND VPWR VPWR _05217_ sky130_fd_sc_hd__a221o_1
Xhold760 data_array.data0\[3\]\[10\] VGND VGND VPWR VPWR net2411 sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 data_array.data1\[13\]\[43\] VGND VGND VPWR VPWR net2422 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold782 data_array.data1\[0\]\[18\] VGND VGND VPWR VPWR net2433 sky130_fd_sc_hd__dlygate4sd3_1
X_11040_ net1751 net1102 net331 VGND VGND VPWR VPWR _02783_ sky130_fd_sc_hd__mux2_1
XFILLER_157_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold793 data_array.data0\[2\]\[59\] VGND VGND VPWR VPWR net2444 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_183_3868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_183_3879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2150 data_array.data1\[12\]\[8\] VGND VGND VPWR VPWR net3801 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2161 data_array.data0\[6\]\[34\] VGND VGND VPWR VPWR net3812 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2172 data_array.data0\[10\]\[7\] VGND VGND VPWR VPWR net3823 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2183 data_array.data1\[13\]\[16\] VGND VGND VPWR VPWR net3834 sky130_fd_sc_hd__dlygate4sd3_1
X_12991_ clknet_leaf_1_clk _01685_ VGND VGND VPWR VPWR data_array.data0\[3\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2194 tag_array.tag1\[6\]\[3\] VGND VGND VPWR VPWR net3845 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1460 data_array.data1\[10\]\[6\] VGND VGND VPWR VPWR net3111 sky130_fd_sc_hd__dlygate4sd3_1
X_11942_ clknet_leaf_222_clk _00750_ VGND VGND VPWR VPWR data_array.data0\[4\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1471 data_array.data0\[14\]\[50\] VGND VGND VPWR VPWR net3122 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1482 data_array.data1\[13\]\[3\] VGND VGND VPWR VPWR net3133 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1493 tag_array.tag1\[13\]\[5\] VGND VGND VPWR VPWR net3144 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_60_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11873_ clknet_leaf_46_clk _00681_ VGND VGND VPWR VPWR data_array.data0\[5\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_13612_ clknet_leaf_218_clk _02241_ VGND VGND VPWR VPWR data_array.data0\[9\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
X_10824_ net1907 net934 net509 VGND VGND VPWR VPWR _02569_ sky130_fd_sc_hd__mux2_1
XFILLER_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13543_ clknet_leaf_123_clk _02172_ VGND VGND VPWR VPWR data_array.data1\[0\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_158_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10755_ net952 net3314 net492 VGND VGND VPWR VPWR _02500_ sky130_fd_sc_hd__mux2_1
XFILLER_9_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_558 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13474_ clknet_leaf_145_clk _02104_ VGND VGND VPWR VPWR tag_array.tag0\[15\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_10686_ net2058 net974 net479 VGND VGND VPWR VPWR _02431_ sky130_fd_sc_hd__mux2_1
XFILLER_173_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12425_ clknet_leaf_47_clk _01119_ VGND VGND VPWR VPWR data_array.data0\[14\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_138_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12356_ clknet_leaf_77_clk _00031_ VGND VGND VPWR VPWR data_array.rdata0\[38\] sky130_fd_sc_hd__dfxtp_1
Xoutput309 net309 VGND VGND VPWR VPWR mem_wdata[51] sky130_fd_sc_hd__buf_2
XFILLER_153_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11307_ net1066 net4548 net800 VGND VGND VPWR VPWR _03050_ sky130_fd_sc_hd__mux2_1
XFILLER_5_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12287_ clknet_leaf_95_clk _01045_ VGND VGND VPWR VPWR tag_array.tag1\[13\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_141_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14026_ clknet_leaf_251_clk _02655_ VGND VGND VPWR VPWR data_array.data1\[6\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_11238_ net1079 net3911 net675 VGND VGND VPWR VPWR _02981_ sky130_fd_sc_hd__mux2_1
XFILLER_150_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_5_27__f_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_5_27__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_171_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11169_ net1099 net2670 net650 VGND VGND VPWR VPWR _02912_ sky130_fd_sc_hd__mux2_1
XFILLER_95_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05730_ net7 fsm.tag_out1\[8\] VGND VGND VPWR VPWR _03247_ sky130_fd_sc_hd__xor2_2
XFILLER_82_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_141_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05661_ net16 fsm.tag_out0\[16\] VGND VGND VPWR VPWR _03178_ sky130_fd_sc_hd__and2b_1
XFILLER_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07400_ data_array.data0\[4\]\[60\] net1411 net1317 data_array.data0\[7\]\[60\] _04644_
+ VGND VGND VPWR VPWR _04645_ sky130_fd_sc_hd__a221o_1
XFILLER_35_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_102_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08380_ net1123 _05489_ VGND VGND VPWR VPWR _05490_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_82_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07331_ data_array.data0\[9\]\[54\] net1547 net1451 data_array.data0\[10\]\[54\]
+ VGND VGND VPWR VPWR _04582_ sky130_fd_sc_hd__a22o_1
X_07262_ net1629 _04513_ _04517_ net1203 VGND VGND VPWR VPWR _04520_ sky130_fd_sc_hd__a22o_1
XFILLER_164_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09001_ net1793 net1020 net419 VGND VGND VPWR VPWR _00756_ sky130_fd_sc_hd__mux2_1
X_06213_ tag_array.tag0\[13\]\[2\] net1559 net1463 tag_array.tag0\[14\]\[2\] VGND
+ VGND VPWR VPWR _03566_ sky130_fd_sc_hd__a22o_1
X_07193_ data_array.data0\[12\]\[41\] net1337 net1243 data_array.data0\[15\]\[41\]
+ _04456_ VGND VGND VPWR VPWR _04457_ sky130_fd_sc_hd__a221o_1
X_06144_ data_array.rdata0\[59\] net1140 net1114 data_array.rdata1\[59\] VGND VGND
+ VPWR VPWR net317 sky130_fd_sc_hd__a22o_1
XFILLER_144_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_148_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_148_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06075_ net1159 net20 fsm.tag_out1\[20\] net1131 VGND VGND VPWR VPWR _03501_ sky130_fd_sc_hd__a22o_1
XFILLER_133_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09903_ net857 net2210 net380 VGND VGND VPWR VPWR _01653_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_165_3532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout503 net504 VGND VGND VPWR VPWR net503 sky130_fd_sc_hd__clkbuf_8
Xfanout514 net515 VGND VGND VPWR VPWR net514 sky130_fd_sc_hd__clkbuf_8
XFILLER_86_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout525 _05599_ VGND VGND VPWR VPWR net525 sky130_fd_sc_hd__clkbuf_4
Xfanout536 net537 VGND VGND VPWR VPWR net536 sky130_fd_sc_hd__buf_2
Xfanout547 _05594_ VGND VGND VPWR VPWR net547 sky130_fd_sc_hd__clkbuf_4
X_09834_ net873 net3344 net390 VGND VGND VPWR VPWR _01585_ sky130_fd_sc_hd__mux2_1
XFILLER_113_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout558 net559 VGND VGND VPWR VPWR net558 sky130_fd_sc_hd__buf_4
XFILLER_112_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout569 net572 VGND VGND VPWR VPWR net569 sky130_fd_sc_hd__buf_2
X_09765_ net1801 net728 net671 VGND VGND VPWR VPWR _01517_ sky130_fd_sc_hd__mux2_1
X_06977_ net1222 _04255_ _04259_ net1173 VGND VGND VPWR VPWR _04261_ sky130_fd_sc_hd__a22o_1
XFILLER_86_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08716_ net1794 net760 net476 VGND VGND VPWR VPWR _00475_ sky130_fd_sc_hd__mux2_1
X_05928_ data_array.rdata1\[32\] net828 net837 VGND VGND VPWR VPWR _03413_ sky130_fd_sc_hd__a21o_1
XFILLER_73_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09696_ net704 net2785 net608 VGND VGND VPWR VPWR _01448_ sky130_fd_sc_hd__mux2_1
XFILLER_132_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08647_ net3182 net735 net506 VGND VGND VPWR VPWR _00406_ sky130_fd_sc_hd__mux2_1
X_05859_ data_array.rdata1\[9\] net832 net841 VGND VGND VPWR VPWR _03367_ sky130_fd_sc_hd__a21o_1
X_08578_ _05595_ net815 VGND VGND VPWR VPWR _05604_ sky130_fd_sc_hd__nand2b_4
XTAP_TAPCELL_ROW_25_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07529_ data_array.data1\[13\]\[8\] net1535 net1439 data_array.data1\[14\]\[8\] VGND
+ VGND VPWR VPWR _04762_ sky130_fd_sc_hd__a22o_1
XFILLER_168_834 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10540_ net1045 net2989 net457 VGND VGND VPWR VPWR _02285_ sky130_fd_sc_hd__mux2_1
XFILLER_41_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10471_ net1061 net2795 net350 VGND VGND VPWR VPWR _02216_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_157_Right_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12210_ clknet_leaf_147_clk _00139_ VGND VGND VPWR VPWR fsm.tag_out0\[17\] sky130_fd_sc_hd__dfxtp_1
X_13190_ clknet_leaf_215_clk _00083_ VGND VGND VPWR VPWR data_array.rdata1\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_157_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12141_ clknet_leaf_143_clk _00949_ VGND VGND VPWR VPWR tag_array.tag0\[12\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_150_222 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12072_ clknet_leaf_46_clk _00880_ VGND VGND VPWR VPWR data_array.data1\[14\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_123_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold590 data_array.data1\[8\]\[24\] VGND VGND VPWR VPWR net2241 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11023_ net1944 net910 net337 VGND VGND VPWR VPWR _02767_ sky130_fd_sc_hd__mux2_1
XFILLER_103_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_86_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12974_ clknet_leaf_169_clk _01668_ VGND VGND VPWR VPWR tag_array.tag0\[4\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_131_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1290 tag_array.tag0\[4\]\[9\] VGND VGND VPWR VPWR net2941 sky130_fd_sc_hd__dlygate4sd3_1
X_11925_ clknet_leaf_226_clk _00733_ VGND VGND VPWR VPWR data_array.data0\[5\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_73_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11856_ clknet_leaf_209_clk _00664_ VGND VGND VPWR VPWR data_array.data0\[7\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10807_ net2191 net1000 net505 VGND VGND VPWR VPWR _02552_ sky130_fd_sc_hd__mux2_1
X_11787_ clknet_leaf_10_clk _00595_ VGND VGND VPWR VPWR data_array.data0\[8\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_159_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13526_ clknet_leaf_200_clk _02155_ VGND VGND VPWR VPWR data_array.data1\[0\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_10738_ net1021 net2936 net492 VGND VGND VPWR VPWR _02483_ sky130_fd_sc_hd__mux2_1
XFILLER_158_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13457_ clknet_leaf_141_clk _02087_ VGND VGND VPWR VPWR tag_array.tag0\[1\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_174_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10669_ net2166 net1040 net478 VGND VGND VPWR VPWR _02414_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_124_Right_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12408_ clknet_leaf_245_clk _01102_ VGND VGND VPWR VPWR data_array.data0\[14\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_126_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13388_ clknet_leaf_19_clk _02018_ VGND VGND VPWR VPWR data_array.data1\[8\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_182_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12339_ clknet_leaf_214_clk _00013_ VGND VGND VPWR VPWR data_array.rdata0\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_141_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2908 data_array.data0\[14\]\[38\] VGND VGND VPWR VPWR net4559 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_101_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2919 data_array.data1\[14\]\[53\] VGND VGND VPWR VPWR net4570 sky130_fd_sc_hd__dlygate4sd3_1
X_06900_ net1176 _04185_ _04189_ net1224 VGND VGND VPWR VPWR _04191_ sky130_fd_sc_hd__a22o_1
X_14009_ clknet_leaf_55_clk _02638_ VGND VGND VPWR VPWR data_array.data1\[5\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
X_07880_ _05080_ _05081_ VGND VGND VPWR VPWR _00096_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_143_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06831_ data_array.data0\[1\]\[8\] net1534 net1438 data_array.data0\[2\]\[8\] VGND
+ VGND VPWR VPWR _04128_ sky130_fd_sc_hd__a22o_1
XFILLER_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_160_3440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09550_ net726 net4520 net620 VGND VGND VPWR VPWR _01303_ sky130_fd_sc_hd__mux2_1
X_06762_ data_array.data0\[4\]\[2\] net1338 net1244 data_array.data0\[7\]\[2\] _04064_
+ VGND VGND VPWR VPWR _04065_ sky130_fd_sc_hd__a221o_1
XFILLER_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08501_ net824 net813 net855 _05556_ VGND VGND VPWR VPWR _05571_ sky130_fd_sc_hd__or4b_4
XTAP_TAPCELL_ROW_121_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_976 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_05713_ _03179_ _03198_ _03204_ _03229_ VGND VGND VPWR VPWR _03230_ sky130_fd_sc_hd__or4_1
X_09481_ net702 net2283 net653 VGND VGND VPWR VPWR _01234_ sky130_fd_sc_hd__mux2_1
X_06693_ tag_array.tag1\[9\]\[21\] net1595 net1499 tag_array.tag1\[10\]\[21\] VGND
+ VGND VPWR VPWR _04002_ sky130_fd_sc_hd__a22o_1
XFILLER_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08432_ net1932 net902 net688 VGND VGND VPWR VPWR _00273_ sky130_fd_sc_hd__mux2_1
X_05644_ net31 fsm.tag_out0\[1\] VGND VGND VPWR VPWR _03161_ sky130_fd_sc_hd__xor2_1
X_08363_ net1908 net992 net691 VGND VGND VPWR VPWR _00250_ sky130_fd_sc_hd__mux2_1
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_158_3391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07314_ data_array.data0\[8\]\[52\] net1357 net1263 data_array.data0\[11\]\[52\]
+ _04566_ VGND VGND VPWR VPWR _04567_ sky130_fd_sc_hd__a221o_1
XFILLER_176_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08294_ net1996 net1084 net686 VGND VGND VPWR VPWR _00227_ sky130_fd_sc_hd__mux2_1
XFILLER_31_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07245_ data_array.data0\[5\]\[46\] net1532 net1436 data_array.data0\[6\]\[46\] VGND
+ VGND VPWR VPWR _04504_ sky130_fd_sc_hd__a22o_1
XFILLER_180_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07176_ _04440_ _04441_ VGND VGND VPWR VPWR _00032_ sky130_fd_sc_hd__or2_1
XFILLER_173_870 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06127_ data_array.rdata0\[42\] net1141 net1115 data_array.rdata1\[42\] VGND VGND
+ VPWR VPWR net299 sky130_fd_sc_hd__a22o_1
XFILLER_11_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06058_ fsm.tag_out0\[11\] net1122 _03492_ VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__a21o_1
XFILLER_160_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1309 net1312 VGND VGND VPWR VPWR net1309 sky130_fd_sc_hd__clkbuf_4
XFILLER_114_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_180_3816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout333 net334 VGND VGND VPWR VPWR net333 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_180_3827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout344 net345 VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__buf_4
Xfanout355 net361 VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__clkbuf_8
Xfanout366 net368 VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__clkbuf_8
XFILLER_59_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout377 _03127_ VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__buf_4
Xclkbuf_5_10__f_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_5_10__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_09817_ net941 net3813 net393 VGND VGND VPWR VPWR _01568_ sky130_fd_sc_hd__mux2_1
XFILLER_143_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout388 net389 VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__buf_4
Xfanout399 net400 VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__buf_4
XFILLER_47_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09748_ net695 net2746 net678 VGND VGND VPWR VPWR _01500_ sky130_fd_sc_hd__mux2_1
XFILLER_43_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09679_ net770 net4507 net606 VGND VGND VPWR VPWR _01431_ sky130_fd_sc_hd__mux2_1
X_11710_ clknet_leaf_164_clk _00518_ VGND VGND VPWR VPWR tag_array.tag0\[9\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_43_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_178_3778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ clknet_leaf_147_clk _01384_ VGND VGND VPWR VPWR tag_array.tag0\[8\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_178_3789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11641_ clknet_leaf_130_clk _00449_ VGND VGND VPWR VPWR tag_array.tag1\[2\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_42_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14360_ clknet_leaf_118_clk _02983_ VGND VGND VPWR VPWR data_array.data1\[10\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11572_ clknet_leaf_132_clk _00380_ VGND VGND VPWR VPWR tag_array.tag1\[5\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13311_ clknet_leaf_125_clk _01941_ VGND VGND VPWR VPWR data_array.data0\[10\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10523_ net1646 net3819 net451 VGND VGND VPWR VPWR _02268_ sky130_fd_sc_hd__mux2_1
Xinput19 cpu_addr[26] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_4
XFILLER_167_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14291_ clknet_leaf_34_clk _02920_ VGND VGND VPWR VPWR data_array.data1\[11\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_109_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13242_ clknet_leaf_64_clk _01872_ VGND VGND VPWR VPWR data_array.data0\[11\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10454_ net353 net3449 net492 VGND VGND VPWR VPWR _02200_ sky130_fd_sc_hd__mux2_1
XFILLER_170_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13173_ clknet_leaf_119_clk _00065_ VGND VGND VPWR VPWR data_array.rdata1\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_184_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10385_ net2039 net352 net635 VGND VGND VPWR VPWR _02131_ sky130_fd_sc_hd__mux2_1
X_12124_ clknet_leaf_180_clk _00932_ VGND VGND VPWR VPWR tag_array.tag0\[12\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12055_ clknet_leaf_263_clk _00863_ VGND VGND VPWR VPWR data_array.data1\[14\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11006_ net1797 net976 net341 VGND VGND VPWR VPWR _02750_ sky130_fd_sc_hd__mux2_1
XFILLER_93_802 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12957_ clknet_leaf_205_clk _01651_ VGND VGND VPWR VPWR data_array.data0\[13\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
X_11908_ clknet_leaf_243_clk _00716_ VGND VGND VPWR VPWR data_array.data0\[5\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12888_ clknet_leaf_13_clk _01582_ VGND VGND VPWR VPWR data_array.data0\[12\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11839_ clknet_leaf_244_clk _00647_ VGND VGND VPWR VPWR data_array.data0\[7\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_16_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13509_ clknet_leaf_268_clk _02138_ VGND VGND VPWR VPWR data_array.data1\[0\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_173_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload202 clknet_leaf_165_clk VGND VGND VPWR VPWR clkload202/Y sky130_fd_sc_hd__clkinvlp_4
X_14489_ clknet_leaf_161_clk _03112_ VGND VGND VPWR VPWR tag_array.dirty0\[8\] sky130_fd_sc_hd__dfxtp_1
Xclkload213 clknet_leaf_109_clk VGND VGND VPWR VPWR clkload213/X sky130_fd_sc_hd__clkbuf_8
X_07030_ data_array.data0\[0\]\[26\] net1339 net1245 data_array.data0\[3\]\[26\] _04308_
+ VGND VGND VPWR VPWR _04309_ sky130_fd_sc_hd__a221o_1
Xclkload224 clknet_leaf_144_clk VGND VGND VPWR VPWR clkload224/X sky130_fd_sc_hd__clkbuf_4
Xclkload235 clknet_leaf_142_clk VGND VGND VPWR VPWR clkload235/Y sky130_fd_sc_hd__clkinv_8
XFILLER_173_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload246 clknet_leaf_147_clk VGND VGND VPWR VPWR clkload246/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_115_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_745 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08981_ net2121 net1102 net420 VGND VGND VPWR VPWR _00736_ sky130_fd_sc_hd__mux2_1
Xhold2705 data_array.data0\[3\]\[53\] VGND VGND VPWR VPWR net4356 sky130_fd_sc_hd__dlygate4sd3_1
X_07932_ data_array.data1\[4\]\[44\] net1398 net1304 data_array.data1\[7\]\[44\] _05128_
+ VGND VGND VPWR VPWR _05129_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_110_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2716 data_array.data1\[3\]\[4\] VGND VGND VPWR VPWR net4367 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2727 data_array.data1\[15\]\[47\] VGND VGND VPWR VPWR net4378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2738 data_array.data1\[6\]\[31\] VGND VGND VPWR VPWR net4389 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2749 data_array.data0\[11\]\[28\] VGND VGND VPWR VPWR net4400 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07863_ data_array.data1\[13\]\[38\] net1588 net1492 data_array.data1\[14\]\[38\]
+ VGND VGND VPWR VPWR _05066_ sky130_fd_sc_hd__a22o_1
XFILLER_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09602_ net941 net3329 net401 VGND VGND VPWR VPWR _01354_ sky130_fd_sc_hd__mux2_1
X_06814_ data_array.data0\[9\]\[7\] net1586 net1490 data_array.data0\[10\]\[7\] VGND
+ VGND VPWR VPWR _04112_ sky130_fd_sc_hd__a22o_1
XFILLER_3_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07794_ data_array.data1\[12\]\[32\] net1330 net1236 data_array.data1\[15\]\[32\]
+ _05002_ VGND VGND VPWR VPWR _05003_ sky130_fd_sc_hd__a221o_1
XFILLER_83_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09533_ net696 net2731 _05567_ VGND VGND VPWR VPWR _01286_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06745_ net1199 _04043_ _04047_ net1625 VGND VGND VPWR VPWR _04050_ sky130_fd_sc_hd__a22o_1
X_09464_ net773 net2479 net658 VGND VGND VPWR VPWR _01217_ sky130_fd_sc_hd__mux2_1
XFILLER_52_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06676_ tag_array.tag1\[12\]\[19\] net1386 net1292 tag_array.tag1\[15\]\[19\] _03986_
+ VGND VGND VPWR VPWR _03987_ sky130_fd_sc_hd__a221o_1
XFILLER_19_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08415_ net140 net75 net1642 VGND VGND VPWR VPWR _05513_ sky130_fd_sc_hd__mux2_1
X_05627_ fsm.state\[2\] _03146_ VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__or2_1
X_09395_ net1087 net3567 net578 VGND VGND VPWR VPWR _01148_ sky130_fd_sc_hd__mux2_1
XFILLER_11_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08346_ net115 net50 net1641 VGND VGND VPWR VPWR _05467_ sky130_fd_sc_hd__mux2_1
XFILLER_178_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_173_3686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08277_ net110 net45 net1638 VGND VGND VPWR VPWR _05421_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_134_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07228_ data_array.data0\[4\]\[44\] net1395 net1301 data_array.data0\[7\]\[44\] _04488_
+ VGND VGND VPWR VPWR _04489_ sky130_fd_sc_hd__a221o_1
XFILLER_137_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07159_ data_array.data0\[13\]\[38\] net1587 net1491 data_array.data0\[14\]\[38\]
+ VGND VGND VPWR VPWR _04426_ sky130_fd_sc_hd__a22o_1
XFILLER_105_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10170_ net867 net3528 net365 VGND VGND VPWR VPWR _01918_ sky130_fd_sc_hd__mux2_1
XFILLER_121_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1106 net1107 VGND VGND VPWR VPWR net1106 sky130_fd_sc_hd__clkbuf_2
XFILLER_121_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1117 net1119 VGND VGND VPWR VPWR net1117 sky130_fd_sc_hd__clkbuf_4
Xfanout1128 net1129 VGND VGND VPWR VPWR net1128 sky130_fd_sc_hd__buf_4
Xfanout1139 net1140 VGND VGND VPWR VPWR net1139 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_802 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13860_ clknet_leaf_234_clk _02489_ VGND VGND VPWR VPWR data_array.data1\[3\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_170_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12811_ clknet_leaf_194_clk _01505_ VGND VGND VPWR VPWR tag_array.tag1\[0\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_13791_ clknet_leaf_200_clk _02420_ VGND VGND VPWR VPWR data_array.data1\[2\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12742_ clknet_leaf_105_clk _01436_ VGND VGND VPWR VPWR tag_array.tag0\[5\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12673_ clknet_leaf_17_clk _01367_ VGND VGND VPWR VPWR data_array.data0\[15\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_190_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_190_clk
+ sky130_fd_sc_hd__clkbuf_8
X_14412_ clknet_leaf_121_clk _03035_ VGND VGND VPWR VPWR data_array.data1\[10\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11624_ clknet_leaf_98_clk _00432_ VGND VGND VPWR VPWR tag_array.tag1\[3\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_13_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14343_ clknet_leaf_192_clk _02972_ VGND VGND VPWR VPWR data_array.data1\[11\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
X_11555_ clknet_leaf_100_clk _00363_ VGND VGND VPWR VPWR tag_array.tag1\[6\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_155_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10506_ net920 net3194 net348 VGND VGND VPWR VPWR _02251_ sky130_fd_sc_hd__mux2_1
XFILLER_144_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14274_ clknet_leaf_203_clk _02903_ VGND VGND VPWR VPWR data_array.data1\[12\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_171_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11486_ clknet_leaf_153_clk _00295_ VGND VGND VPWR VPWR tag_array.valid0\[0\] sky130_fd_sc_hd__dfxtp_1
X_13225_ clknet_leaf_119_clk _00122_ VGND VGND VPWR VPWR data_array.rdata1\[62\] sky130_fd_sc_hd__dfxtp_1
X_10437_ net2826 net907 net661 VGND VGND VPWR VPWR _02183_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_78_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13156_ clknet_leaf_187_clk _01850_ VGND VGND VPWR VPWR tag_array.tag1\[8\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_10368_ net727 net2717 net539 VGND VGND VPWR VPWR _02115_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12107_ clknet_leaf_5_clk _00915_ VGND VGND VPWR VPWR data_array.data1\[14\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13087_ clknet_leaf_77_clk _01781_ VGND VGND VPWR VPWR data_array.data1\[13\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_72_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10299_ net2373 net966 net640 VGND VGND VPWR VPWR _02046_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1640 net1641 VGND VGND VPWR VPWR net1640 sky130_fd_sc_hd__buf_4
X_12038_ clknet_leaf_40_clk _00846_ VGND VGND VPWR VPWR data_array.data0\[6\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout1651 net163 VGND VGND VPWR VPWR net1651 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13989_ clknet_leaf_39_clk _02618_ VGND VGND VPWR VPWR data_array.data1\[5\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_87_Right_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06530_ tag_array.tag1\[1\]\[6\] net1552 net1456 tag_array.tag1\[2\]\[6\] VGND VGND
+ VPWR VPWR _03854_ sky130_fd_sc_hd__a22o_1
XFILLER_92_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06461_ _03790_ _03791_ VGND VGND VPWR VPWR _00147_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_138_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_181_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_181_clk
+ sky130_fd_sc_hd__clkbuf_8
X_08200_ _03136_ _03147_ VGND VGND VPWR VPWR _05368_ sky130_fd_sc_hd__nor2_1
XFILLER_166_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09180_ net758 net2762 net629 VGND VGND VPWR VPWR _00934_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_155_3350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06392_ tag_array.tag0\[4\]\[18\] net1407 net1313 tag_array.tag0\[7\]\[18\] _03728_
+ VGND VGND VPWR VPWR _03729_ sky130_fd_sc_hd__a221o_1
XFILLER_175_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08131_ net1635 _05303_ _05307_ net1209 VGND VGND VPWR VPWR _05310_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_79_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08062_ data_array.data1\[8\]\[56\] net1341 net1247 data_array.data1\[11\]\[56\]
+ _05246_ VGND VGND VPWR VPWR _05247_ sky130_fd_sc_hd__a221o_1
XFILLER_107_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07013_ data_array.data0\[12\]\[25\] net1329 net1235 data_array.data0\[15\]\[25\]
+ _04292_ VGND VGND VPWR VPWR _04293_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_96_Right_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2502 tag_array.tag0\[1\]\[20\] VGND VGND VPWR VPWR net4153 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_142_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2513 data_array.data0\[7\]\[21\] VGND VGND VPWR VPWR net4164 sky130_fd_sc_hd__dlygate4sd3_1
X_08964_ net910 net2766 net427 VGND VGND VPWR VPWR _00720_ sky130_fd_sc_hd__mux2_1
XFILLER_103_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2524 data_array.data0\[14\]\[22\] VGND VGND VPWR VPWR net4175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2535 data_array.data1\[11\]\[21\] VGND VGND VPWR VPWR net4186 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1801 data_array.data0\[14\]\[15\] VGND VGND VPWR VPWR net3452 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2546 data_array.data0\[10\]\[41\] VGND VGND VPWR VPWR net4197 sky130_fd_sc_hd__dlygate4sd3_1
X_07915_ data_array.data1\[8\]\[43\] net1378 net1284 data_array.data1\[11\]\[43\]
+ _05112_ VGND VGND VPWR VPWR _05113_ sky130_fd_sc_hd__a221o_1
Xhold1812 data_array.data0\[5\]\[60\] VGND VGND VPWR VPWR net3463 sky130_fd_sc_hd__dlygate4sd3_1
X_08895_ net927 net3927 net434 VGND VGND VPWR VPWR _00652_ sky130_fd_sc_hd__mux2_1
Xhold2557 tag_array.tag1\[3\]\[14\] VGND VGND VPWR VPWR net4208 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2568 data_array.data0\[11\]\[25\] VGND VGND VPWR VPWR net4219 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1823 data_array.data0\[6\]\[23\] VGND VGND VPWR VPWR net3474 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2579 data_array.data0\[7\]\[55\] VGND VGND VPWR VPWR net4230 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1834 tag_array.tag0\[8\]\[10\] VGND VGND VPWR VPWR net3485 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1845 data_array.data0\[11\]\[6\] VGND VGND VPWR VPWR net3496 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_25_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07846_ net1186 _05045_ _05049_ net1231 VGND VGND VPWR VPWR _05051_ sky130_fd_sc_hd__a22o_1
XFILLER_151_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1856 tag_array.tag0\[9\]\[15\] VGND VGND VPWR VPWR net3507 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_110_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1867 tag_array.tag1\[7\]\[0\] VGND VGND VPWR VPWR net3518 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1878 data_array.data1\[5\]\[20\] VGND VGND VPWR VPWR net3529 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1889 data_array.data1\[15\]\[43\] VGND VGND VPWR VPWR net3540 sky130_fd_sc_hd__dlygate4sd3_1
X_07777_ data_array.data1\[1\]\[30\] net1583 net1487 data_array.data1\[2\]\[30\] VGND
+ VGND VPWR VPWR _04988_ sky130_fd_sc_hd__a22o_1
XFILLER_140_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06728_ tag_array.tag1\[5\]\[24\] net1562 net1466 tag_array.tag1\[6\]\[24\] VGND
+ VGND VPWR VPWR _04034_ sky130_fd_sc_hd__a22o_1
X_09516_ net762 net3991 net623 VGND VGND VPWR VPWR _01269_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_175_3715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_175_3726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09447_ net879 net3137 net582 VGND VGND VPWR VPWR _01200_ sky130_fd_sc_hd__mux2_1
X_06659_ _03970_ _03971_ VGND VGND VPWR VPWR _00164_ sky130_fd_sc_hd__or2_1
XFILLER_24_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_172_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_172_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_33_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_12 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09378_ net889 net4286 net403 VGND VGND VPWR VPWR _01131_ sky130_fd_sc_hd__mux2_1
XFILLER_40_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08329_ net1128 _05455_ VGND VGND VPWR VPWR _05456_ sky130_fd_sc_hd__and2_1
XFILLER_32_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11340_ net934 net3841 net802 VGND VGND VPWR VPWR _03083_ sky130_fd_sc_hd__mux2_1
X_11271_ net945 net4406 net673 VGND VGND VPWR VPWR _03014_ sky130_fd_sc_hd__mux2_1
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13010_ clknet_leaf_268_clk _01704_ VGND VGND VPWR VPWR data_array.data0\[3\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_37_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10222_ net916 net4255 net359 VGND VGND VPWR VPWR _01969_ sky130_fd_sc_hd__mux2_1
XFILLER_140_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_5_8__f_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_5_8__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_10153_ net933 net4497 net368 VGND VGND VPWR VPWR _01901_ sky130_fd_sc_hd__mux2_1
XFILLER_58_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10084_ net2172 net786 net635 VGND VGND VPWR VPWR _01833_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13912_ clknet_leaf_212_clk _02541_ VGND VGND VPWR VPWR data_array.data1\[4\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_114_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13843_ clknet_leaf_35_clk _02472_ VGND VGND VPWR VPWR data_array.data1\[3\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_18_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13774_ clknet_leaf_268_clk _02403_ VGND VGND VPWR VPWR data_array.data1\[2\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_10986_ net1819 net1058 net338 VGND VGND VPWR VPWR _02730_ sky130_fd_sc_hd__mux2_1
X_12725_ clknet_leaf_153_clk _01419_ VGND VGND VPWR VPWR tag_array.tag0\[7\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_163_clk clknet_5_25__leaf_clk VGND VGND VPWR VPWR clknet_leaf_163_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12656_ clknet_leaf_73_clk _01350_ VGND VGND VPWR VPWR data_array.data0\[15\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_175_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11607_ clknet_leaf_129_clk _00415_ VGND VGND VPWR VPWR tag_array.tag1\[4\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_96_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12587_ clknet_leaf_161_clk _01281_ VGND VGND VPWR VPWR tag_array.tag0\[10\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14326_ clknet_leaf_244_clk _02955_ VGND VGND VPWR VPWR data_array.data1\[11\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
X_11538_ clknet_leaf_193_clk _00346_ VGND VGND VPWR VPWR tag_array.tag1\[6\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_171_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_423 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold408 data_array.data1\[1\]\[57\] VGND VGND VPWR VPWR net2059 sky130_fd_sc_hd__dlygate4sd3_1
Xhold419 data_array.data0\[1\]\[47\] VGND VGND VPWR VPWR net2070 sky130_fd_sc_hd__dlygate4sd3_1
X_11469_ clknet_leaf_207_clk _00279_ VGND VGND VPWR VPWR data_array.data0\[0\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
X_14257_ clknet_leaf_258_clk _02886_ VGND VGND VPWR VPWR data_array.data1\[12\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_74_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1022 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13208_ clknet_leaf_14_clk _00103_ VGND VGND VPWR VPWR data_array.rdata1\[45\] sky130_fd_sc_hd__dfxtp_1
X_14188_ clknet_leaf_85_clk _02817_ VGND VGND VPWR VPWR data_array.data0\[2\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_112_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13139_ clknet_leaf_232_clk _01833_ VGND VGND VPWR VPWR tag_array.tag1\[8\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_98_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05961_ data_array.rdata1\[43\] net833 net842 VGND VGND VPWR VPWR _03435_ sky130_fd_sc_hd__a21o_1
Xhold1108 data_array.data1\[6\]\[29\] VGND VGND VPWR VPWR net2759 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1119 data_array.data1\[9\]\[46\] VGND VGND VPWR VPWR net2770 sky130_fd_sc_hd__dlygate4sd3_1
X_07700_ data_array.data1\[5\]\[23\] net1550 net1454 data_array.data1\[6\]\[23\] VGND
+ VGND VPWR VPWR _04918_ sky130_fd_sc_hd__a22o_1
Xfanout1470 net1518 VGND VGND VPWR VPWR net1470 sky130_fd_sc_hd__buf_2
X_08680_ net702 net3484 net493 VGND VGND VPWR VPWR _00439_ sky130_fd_sc_hd__mux2_1
Xfanout1481 net1483 VGND VGND VPWR VPWR net1481 sky130_fd_sc_hd__clkbuf_4
X_05892_ data_array.rdata1\[20\] net834 net843 VGND VGND VPWR VPWR _03389_ sky130_fd_sc_hd__a21o_1
XFILLER_94_963 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1492 net1494 VGND VGND VPWR VPWR net1492 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07631_ data_array.data1\[0\]\[17\] net1336 net1242 data_array.data1\[3\]\[17\] _04854_
+ VGND VGND VPWR VPWR _04855_ sky130_fd_sc_hd__a221o_1
XFILLER_19_592 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07562_ data_array.data1\[9\]\[11\] net1574 net1478 data_array.data1\[10\]\[11\]
+ VGND VGND VPWR VPWR _04792_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_105_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09301_ net774 net2642 net546 VGND VGND VPWR VPWR _01055_ sky130_fd_sc_hd__mux2_1
X_06513_ tag_array.tag1\[4\]\[4\] net1362 net1268 tag_array.tag1\[7\]\[4\] _03838_
+ VGND VGND VPWR VPWR _03839_ sky130_fd_sc_hd__a221o_1
X_07493_ net1630 _04723_ _04727_ net1204 VGND VGND VPWR VPWR _04730_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_154_clk clknet_5_28__leaf_clk VGND VGND VPWR VPWR clknet_leaf_154_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_181_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09232_ net752 net3464 net646 VGND VGND VPWR VPWR _00986_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_153_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06444_ tag_array.tag0\[13\]\[23\] net1598 net1502 tag_array.tag0\[14\]\[23\] VGND
+ VGND VPWR VPWR _03776_ sky130_fd_sc_hd__a22o_1
XFILLER_21_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_170_3623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09163_ net890 net3677 net568 VGND VGND VPWR VPWR _00917_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_170_3634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06375_ tag_array.tag0\[12\]\[17\] net1405 net1311 tag_array.tag0\[15\]\[17\] _03712_
+ VGND VGND VPWR VPWR _03713_ sky130_fd_sc_hd__a221o_1
X_08114_ data_array.data1\[1\]\[61\] net1550 net1454 data_array.data1\[2\]\[61\] VGND
+ VGND VPWR VPWR _05294_ sky130_fd_sc_hd__a22o_1
X_09094_ net909 net3838 net411 VGND VGND VPWR VPWR _00848_ sky130_fd_sc_hd__mux2_1
XFILLER_174_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08045_ _05230_ _05231_ VGND VGND VPWR VPWR _00113_ sky130_fd_sc_hd__or2_1
Xhold920 data_array.data1\[2\]\[56\] VGND VGND VPWR VPWR net2571 sky130_fd_sc_hd__dlygate4sd3_1
Xhold931 tag_array.tag0\[3\]\[10\] VGND VGND VPWR VPWR net2582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold942 data_array.data0\[4\]\[13\] VGND VGND VPWR VPWR net2593 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold953 data_array.data1\[13\]\[27\] VGND VGND VPWR VPWR net2604 sky130_fd_sc_hd__dlygate4sd3_1
Xhold964 data_array.data0\[9\]\[2\] VGND VGND VPWR VPWR net2615 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold975 data_array.data0\[8\]\[34\] VGND VGND VPWR VPWR net2626 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold986 tag_array.tag1\[13\]\[18\] VGND VGND VPWR VPWR net2637 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_168_3585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold997 tag_array.tag1\[4\]\[24\] VGND VGND VPWR VPWR net2648 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_168_3596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09996_ net1100 net2627 net555 VGND VGND VPWR VPWR _01745_ sky130_fd_sc_hd__mux2_1
Xhold2310 tag_array.tag0\[8\]\[11\] VGND VGND VPWR VPWR net3961 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_134_Left_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2321 data_array.data1\[14\]\[34\] VGND VGND VPWR VPWR net3972 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2332 data_array.data0\[11\]\[53\] VGND VGND VPWR VPWR net3983 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2343 data_array.data0\[14\]\[23\] VGND VGND VPWR VPWR net3994 sky130_fd_sc_hd__dlygate4sd3_1
X_08947_ net976 net4357 net430 VGND VGND VPWR VPWR _00703_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2354 data_array.data0\[7\]\[31\] VGND VGND VPWR VPWR net4005 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1620 data_array.data1\[10\]\[61\] VGND VGND VPWR VPWR net3271 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2365 tag_array.tag0\[1\]\[19\] VGND VGND VPWR VPWR net4016 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2376 tag_array.tag1\[13\]\[15\] VGND VGND VPWR VPWR net4027 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1631 data_array.data0\[5\]\[12\] VGND VGND VPWR VPWR net3282 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1642 tag_array.tag1\[7\]\[10\] VGND VGND VPWR VPWR net3293 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2387 tag_array.tag0\[3\]\[5\] VGND VGND VPWR VPWR net4038 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2398 tag_array.dirty1\[15\] VGND VGND VPWR VPWR net4049 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1653 data_array.data1\[3\]\[43\] VGND VGND VPWR VPWR net3304 sky130_fd_sc_hd__dlygate4sd3_1
X_08878_ net992 net4044 net438 VGND VGND VPWR VPWR _00635_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1664 tag_array.tag0\[5\]\[18\] VGND VGND VPWR VPWR net3315 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1675 tag_array.tag0\[10\]\[13\] VGND VGND VPWR VPWR net3326 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1686 data_array.data0\[3\]\[52\] VGND VGND VPWR VPWR net3337 sky130_fd_sc_hd__dlygate4sd3_1
X_07829_ data_array.data1\[4\]\[35\] net1335 net1241 data_array.data1\[7\]\[35\] _05034_
+ VGND VGND VPWR VPWR _05035_ sky130_fd_sc_hd__a221o_1
Xhold1697 tag_array.tag1\[14\]\[8\] VGND VGND VPWR VPWR net3348 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10840_ net2139 net870 net510 VGND VGND VPWR VPWR _02585_ sky130_fd_sc_hd__mux2_1
XFILLER_71_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10771_ net890 net3563 net492 VGND VGND VPWR VPWR _02516_ sky130_fd_sc_hd__mux2_1
XFILLER_40_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_145_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_145_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_143_Left_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12510_ clknet_leaf_121_clk _01204_ VGND VGND VPWR VPWR data_array.data1\[9\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
X_13490_ clknet_leaf_155_clk _02120_ VGND VGND VPWR VPWR tag_array.tag0\[15\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_139_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12441_ clknet_leaf_51_clk _01135_ VGND VGND VPWR VPWR data_array.data0\[14\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12372_ clknet_leaf_214_clk _00049_ VGND VGND VPWR VPWR data_array.rdata0\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_176_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11323_ net1000 net3361 net798 VGND VGND VPWR VPWR _03066_ sky130_fd_sc_hd__mux2_1
X_14111_ clknet_leaf_225_clk _02740_ VGND VGND VPWR VPWR data_array.data0\[1\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_4_0_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_0_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14042_ clknet_leaf_18_clk _02671_ VGND VGND VPWR VPWR data_array.data1\[6\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_109_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11254_ net1014 net4440 net681 VGND VGND VPWR VPWR _02997_ sky130_fd_sc_hd__mux2_1
XFILLER_122_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_152_Left_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10205_ net986 net3431 net358 VGND VGND VPWR VPWR _01952_ sky130_fd_sc_hd__mux2_1
XFILLER_140_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_843 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11185_ net1035 net4171 net656 VGND VGND VPWR VPWR _02928_ sky130_fd_sc_hd__mux2_1
XFILLER_121_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10136_ net1003 net4203 net365 VGND VGND VPWR VPWR _01884_ sky130_fd_sc_hd__mux2_1
XFILLER_95_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10067_ net754 net3747 net600 VGND VGND VPWR VPWR _01816_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_89_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_996 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13826_ clknet_leaf_202_clk _02455_ VGND VGND VPWR VPWR data_array.data1\[2\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_91_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_161_Left_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_136_clk clknet_5_31__leaf_clk VGND VGND VPWR VPWR clknet_leaf_136_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13757_ clknet_leaf_7_clk _02386_ VGND VGND VPWR VPWR data_array.data1\[1\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
X_10969_ net864 net4565 net529 VGND VGND VPWR VPWR _02714_ sky130_fd_sc_hd__mux2_1
X_12708_ clknet_leaf_164_clk _01402_ VGND VGND VPWR VPWR tag_array.tag0\[7\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13688_ clknet_leaf_75_clk _02317_ VGND VGND VPWR VPWR data_array.data1\[15\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_148_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12639_ clknet_leaf_226_clk _01333_ VGND VGND VPWR VPWR data_array.data0\[15\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_157_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06160_ tag_array.valid0\[8\] net1407 net1313 tag_array.valid0\[11\] _03512_ VGND
+ VGND VPWR VPWR _03517_ sky130_fd_sc_hd__a221o_1
XFILLER_156_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_935 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_732 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold205 data_array.data0\[8\]\[31\] VGND VGND VPWR VPWR net1856 sky130_fd_sc_hd__dlygate4sd3_1
X_14309_ clknet_leaf_40_clk _02938_ VGND VGND VPWR VPWR data_array.data1\[11\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_06091_ data_array.rdata0\[6\] net1134 net1112 data_array.rdata1\[6\] VGND VGND VPWR
+ VPWR net323 sky130_fd_sc_hd__a22o_1
Xhold216 tag_array.tag1\[2\]\[1\] VGND VGND VPWR VPWR net1867 sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 data_array.data0\[8\]\[8\] VGND VGND VPWR VPWR net1878 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_170_Left_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold238 data_array.data0\[2\]\[37\] VGND VGND VPWR VPWR net1889 sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 data_array.data1\[4\]\[50\] VGND VGND VPWR VPWR net1900 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout707 _05407_ VGND VGND VPWR VPWR net707 sky130_fd_sc_hd__dlymetal6s2s_1
X_09850_ net1069 net2643 net384 VGND VGND VPWR VPWR _01600_ sky130_fd_sc_hd__mux2_1
Xfanout718 net721 VGND VGND VPWR VPWR net718 sky130_fd_sc_hd__clkbuf_2
Xfanout729 _05397_ VGND VGND VPWR VPWR net729 sky130_fd_sc_hd__clkbuf_2
XFILLER_98_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08801_ net2150 net1043 net442 VGND VGND VPWR VPWR _00559_ sky130_fd_sc_hd__mux2_1
X_09781_ net1085 net2508 net386 VGND VGND VPWR VPWR _01532_ sky130_fd_sc_hd__mux2_1
X_06993_ data_array.data0\[0\]\[23\] net1366 net1272 data_array.data0\[3\]\[23\] _04274_
+ VGND VGND VPWR VPWR _04275_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_146_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05944_ net129 net1152 _03422_ _03423_ VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__a22o_1
X_08732_ net2828 net694 net470 VGND VGND VPWR VPWR _00491_ sky130_fd_sc_hd__mux2_1
XFILLER_22_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_163_3493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08663_ net772 net2953 net500 VGND VGND VPWR VPWR _00422_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05875_ net104 net1156 _03376_ _03377_ VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__a22o_1
XFILLER_81_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07614_ net1632 _04833_ _04837_ net1206 VGND VGND VPWR VPWR _04840_ sky130_fd_sc_hd__a22o_1
X_08594_ net746 net3672 net534 VGND VGND VPWR VPWR _00353_ sky130_fd_sc_hd__mux2_1
XFILLER_53_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07545_ data_array.data1\[12\]\[9\] net1391 net1297 data_array.data1\[15\]\[9\] _04776_
+ VGND VGND VPWR VPWR _04777_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_127_clk clknet_5_30__leaf_clk VGND VGND VPWR VPWR clknet_leaf_127_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_138_Right_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07476_ data_array.data1\[5\]\[3\] net1540 net1444 data_array.data1\[6\]\[3\] VGND
+ VGND VPWR VPWR _04714_ sky130_fd_sc_hd__a22o_1
XFILLER_22_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09215_ net720 net4247 net630 VGND VGND VPWR VPWR _00969_ sky130_fd_sc_hd__mux2_1
X_06427_ net1182 _03755_ _03759_ net1234 VGND VGND VPWR VPWR _03761_ sky130_fd_sc_hd__a22o_1
XFILLER_10_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09146_ net959 net4543 net574 VGND VGND VPWR VPWR _00900_ sky130_fd_sc_hd__mux2_1
X_06358_ tag_array.tag0\[5\]\[15\] net1593 net1497 tag_array.tag0\[6\]\[15\] VGND
+ VGND VPWR VPWR _03698_ sky130_fd_sc_hd__a22o_1
XFILLER_5_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09077_ net976 net4145 net414 VGND VGND VPWR VPWR _00831_ sky130_fd_sc_hd__mux2_1
X_06289_ tag_array.tag0\[0\]\[9\] net1409 net1315 tag_array.tag0\[3\]\[9\] _03634_
+ VGND VGND VPWR VPWR _03635_ sky130_fd_sc_hd__a221o_1
XFILLER_107_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08028_ data_array.data1\[13\]\[53\] net1523 net1427 data_array.data1\[14\]\[53\]
+ VGND VGND VPWR VPWR _05216_ sky130_fd_sc_hd__a22o_1
XFILLER_100_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold750 data_array.data1\[10\]\[60\] VGND VGND VPWR VPWR net2401 sky130_fd_sc_hd__dlygate4sd3_1
Xhold761 data_array.data1\[1\]\[52\] VGND VGND VPWR VPWR net2412 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold772 data_array.data1\[9\]\[34\] VGND VGND VPWR VPWR net2423 sky130_fd_sc_hd__dlygate4sd3_1
Xhold783 data_array.data1\[9\]\[13\] VGND VGND VPWR VPWR net2434 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold794 data_array.data0\[2\]\[27\] VGND VGND VPWR VPWR net2445 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_183_3869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_34 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09979_ net912 net4229 net375 VGND VGND VPWR VPWR _01728_ sky130_fd_sc_hd__mux2_1
Xhold2140 data_array.data1\[6\]\[58\] VGND VGND VPWR VPWR net3791 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2151 data_array.data1\[14\]\[31\] VGND VGND VPWR VPWR net3802 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2162 data_array.data0\[12\]\[42\] VGND VGND VPWR VPWR net3813 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2173 data_array.data1\[7\]\[0\] VGND VGND VPWR VPWR net3824 sky130_fd_sc_hd__dlygate4sd3_1
X_12990_ clknet_leaf_210_clk _01684_ VGND VGND VPWR VPWR data_array.data0\[3\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2184 tag_array.tag0\[3\]\[4\] VGND VGND VPWR VPWR net3835 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1450 data_array.data1\[14\]\[61\] VGND VGND VPWR VPWR net3101 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2195 data_array.data0\[7\]\[0\] VGND VGND VPWR VPWR net3846 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1461 tag_array.tag1\[3\]\[23\] VGND VGND VPWR VPWR net3112 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11941_ clknet_leaf_63_clk _00749_ VGND VGND VPWR VPWR data_array.data0\[4\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1472 data_array.data0\[6\]\[61\] VGND VGND VPWR VPWR net3123 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1483 tag_array.tag0\[0\]\[9\] VGND VGND VPWR VPWR net3134 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1494 tag_array.tag0\[2\]\[8\] VGND VGND VPWR VPWR net3145 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11872_ clknet_leaf_112_clk _00680_ VGND VGND VPWR VPWR data_array.data0\[5\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_13611_ clknet_leaf_114_clk _02240_ VGND VGND VPWR VPWR data_array.data0\[9\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
X_10823_ net1744 net937 net507 VGND VGND VPWR VPWR _02568_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_118_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_118_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_105_Right_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13542_ clknet_leaf_240_clk _02171_ VGND VGND VPWR VPWR data_array.data1\[0\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
X_10754_ net958 net3139 net498 VGND VGND VPWR VPWR _02499_ sky130_fd_sc_hd__mux2_1
X_10685_ net4368 net977 net484 VGND VGND VPWR VPWR _02430_ sky130_fd_sc_hd__mux2_1
XFILLER_9_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13473_ clknet_leaf_181_clk _02103_ VGND VGND VPWR VPWR tag_array.tag0\[15\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_12424_ clknet_leaf_93_clk _01118_ VGND VGND VPWR VPWR data_array.data0\[14\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_139_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12355_ clknet_leaf_214_clk _00030_ VGND VGND VPWR VPWR data_array.rdata0\[37\] sky130_fd_sc_hd__dfxtp_1
X_11306_ net1071 net3453 net804 VGND VGND VPWR VPWR _03049_ sky130_fd_sc_hd__mux2_1
X_12286_ clknet_leaf_187_clk _01044_ VGND VGND VPWR VPWR tag_array.tag1\[13\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_107_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11237_ net1082 net4101 net682 VGND VGND VPWR VPWR _02980_ sky130_fd_sc_hd__mux2_1
X_14025_ clknet_leaf_267_clk _02654_ VGND VGND VPWR VPWR data_array.data1\[6\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_11168_ net1101 net4545 net649 VGND VGND VPWR VPWR _02911_ sky130_fd_sc_hd__mux2_1
XFILLER_45_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10119_ net1069 net3301 net368 VGND VGND VPWR VPWR _01867_ sky130_fd_sc_hd__mux2_1
X_11099_ net2265 net866 net330 VGND VGND VPWR VPWR _02842_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_69_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_141_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05660_ _03162_ _03166_ _03171_ _03176_ VGND VGND VPWR VPWR _03177_ sky130_fd_sc_hd__or4_4
XFILLER_91_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13809_ clknet_leaf_257_clk _02438_ VGND VGND VPWR VPWR data_array.data1\[2\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_109_clk clknet_5_27__leaf_clk VGND VGND VPWR VPWR clknet_leaf_109_clk
+ sky130_fd_sc_hd__clkbuf_8
X_07330_ _04580_ _04581_ VGND VGND VPWR VPWR _00048_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_82_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07261_ data_array.data0\[0\]\[47\] net1387 net1293 data_array.data0\[3\]\[47\] _04518_
+ VGND VGND VPWR VPWR _04519_ sky130_fd_sc_hd__a221o_1
X_09000_ net2580 net1026 net421 VGND VGND VPWR VPWR _00755_ sky130_fd_sc_hd__mux2_1
X_06212_ tag_array.tag0\[4\]\[2\] net1370 net1276 tag_array.tag0\[7\]\[2\] _03564_
+ VGND VGND VPWR VPWR _03565_ sky130_fd_sc_hd__a221o_1
X_07192_ data_array.data0\[13\]\[41\] net1527 net1431 data_array.data0\[14\]\[41\]
+ VGND VGND VPWR VPWR _04456_ sky130_fd_sc_hd__a22o_1
X_06143_ data_array.rdata0\[58\] net1136 net1117 data_array.rdata1\[58\] VGND VGND
+ VPWR VPWR net316 sky130_fd_sc_hd__a22o_1
XFILLER_144_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06074_ fsm.tag_out0\[19\] net1121 _03500_ VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_148_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09902_ net861 net2813 net385 VGND VGND VPWR VPWR _01652_ sky130_fd_sc_hd__mux2_1
XFILLER_99_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout504 net513 VGND VGND VPWR VPWR net504 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_165_3533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout515 net518 VGND VGND VPWR VPWR net515 sky130_fd_sc_hd__clkbuf_8
Xfanout526 net527 VGND VGND VPWR VPWR net526 sky130_fd_sc_hd__clkbuf_8
X_09833_ net877 net4306 net389 VGND VGND VPWR VPWR _01584_ sky130_fd_sc_hd__mux2_1
Xfanout537 _05598_ VGND VGND VPWR VPWR net537 sky130_fd_sc_hd__clkbuf_4
XFILLER_113_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout548 net553 VGND VGND VPWR VPWR net548 sky130_fd_sc_hd__buf_4
Xfanout559 net560 VGND VGND VPWR VPWR net559 sky130_fd_sc_hd__buf_4
XFILLER_100_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09764_ net1890 net730 net670 VGND VGND VPWR VPWR _01516_ sky130_fd_sc_hd__mux2_1
X_06976_ net1621 _04253_ _04257_ net1195 VGND VGND VPWR VPWR _04260_ sky130_fd_sc_hd__a22o_1
XFILLER_132_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08715_ net2764 net764 net475 VGND VGND VPWR VPWR _00474_ sky130_fd_sc_hd__mux2_1
X_05927_ data_array.rdata0\[32\] net846 net1142 VGND VGND VPWR VPWR _03412_ sky130_fd_sc_hd__o21a_1
XFILLER_6_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09695_ net709 net4030 net607 VGND VGND VPWR VPWR _01447_ sky130_fd_sc_hd__mux2_1
XFILLER_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08646_ net1771 net740 net511 VGND VGND VPWR VPWR _00405_ sky130_fd_sc_hd__mux2_1
X_05858_ data_array.rdata0\[9\] net850 net1147 VGND VGND VPWR VPWR _03366_ sky130_fd_sc_hd__o21a_1
XFILLER_81_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08577_ net1723 net470 VGND VGND VPWR VPWR _00339_ sky130_fd_sc_hd__or2_1
X_05789_ _03251_ _03258_ _03270_ _03278_ VGND VGND VPWR VPWR _03306_ sky130_fd_sc_hd__or4_1
XFILLER_23_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07528_ _04760_ _04761_ VGND VGND VPWR VPWR _00125_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_25_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07459_ data_array.data1\[4\]\[1\] net1330 net1236 data_array.data1\[7\]\[1\] _04698_
+ VGND VGND VPWR VPWR _04699_ sky130_fd_sc_hd__a221o_1
X_10470_ net1065 net2556 net348 VGND VGND VPWR VPWR _02215_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09129_ net1024 net3398 net567 VGND VGND VPWR VPWR _00883_ sky130_fd_sc_hd__mux2_1
XFILLER_108_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12140_ clknet_leaf_182_clk _00948_ VGND VGND VPWR VPWR tag_array.tag0\[12\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12071_ clknet_leaf_250_clk _00879_ VGND VGND VPWR VPWR data_array.data1\[14\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold580 data_array.data1\[4\]\[49\] VGND VGND VPWR VPWR net2231 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_173_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold591 data_array.data0\[8\]\[30\] VGND VGND VPWR VPWR net2242 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11022_ net1739 net912 net341 VGND VGND VPWR VPWR _02766_ sky130_fd_sc_hd__mux2_1
XFILLER_1_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12973_ clknet_leaf_139_clk _01667_ VGND VGND VPWR VPWR tag_array.tag0\[4\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1280 data_array.data0\[9\]\[17\] VGND VGND VPWR VPWR net2931 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1291 data_array.data0\[5\]\[3\] VGND VGND VPWR VPWR net2942 sky130_fd_sc_hd__dlygate4sd3_1
X_11924_ clknet_leaf_109_clk _00732_ VGND VGND VPWR VPWR data_array.data0\[5\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_45_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11855_ clknet_leaf_236_clk _00663_ VGND VGND VPWR VPWR data_array.data0\[7\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_64_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10806_ net1843 net1004 net504 VGND VGND VPWR VPWR _02551_ sky130_fd_sc_hd__mux2_1
X_11786_ clknet_leaf_207_clk _00594_ VGND VGND VPWR VPWR data_array.data0\[8\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_41_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13525_ clknet_leaf_24_clk _02154_ VGND VGND VPWR VPWR data_array.data1\[0\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_41_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10737_ net1025 net3579 net494 VGND VGND VPWR VPWR _02482_ sky130_fd_sc_hd__mux2_1
X_13456_ clknet_leaf_163_clk _02086_ VGND VGND VPWR VPWR tag_array.tag0\[1\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_139_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10668_ net2398 net1044 net481 VGND VGND VPWR VPWR _02413_ sky130_fd_sc_hd__mux2_1
XFILLER_12_1024 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12407_ clknet_leaf_262_clk _01101_ VGND VGND VPWR VPWR data_array.data0\[14\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_13387_ clknet_leaf_118_clk _02017_ VGND VGND VPWR VPWR data_array.data1\[8\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_10599_ net2035 net1067 net471 VGND VGND VPWR VPWR _02344_ sky130_fd_sc_hd__mux2_1
XFILLER_127_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12338_ clknet_leaf_131_clk _00012_ VGND VGND VPWR VPWR data_array.rdata0\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12269_ clknet_leaf_167_clk _01027_ VGND VGND VPWR VPWR tag_array.tag1\[13\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2909 data_array.data0\[6\]\[32\] VGND VGND VPWR VPWR net4560 sky130_fd_sc_hd__dlygate4sd3_1
X_14008_ clknet_leaf_71_clk _02637_ VGND VGND VPWR VPWR data_array.data1\[5\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_143_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06830_ data_array.data0\[8\]\[8\] net1343 net1249 data_array.data0\[11\]\[8\] _04126_
+ VGND VGND VPWR VPWR _04127_ sky130_fd_sc_hd__a221o_1
XFILLER_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_3430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06761_ data_array.data0\[5\]\[2\] net1529 net1433 data_array.data0\[6\]\[2\] VGND
+ VGND VPWR VPWR _04064_ sky130_fd_sc_hd__a22o_1
XFILLER_37_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08500_ _03507_ _03514_ net825 VGND VGND VPWR VPWR _05570_ sky130_fd_sc_hd__or3_1
X_05712_ fsm.tag_out0\[2\] net32 VGND VGND VPWR VPWR _03229_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_121_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06692_ _04000_ _04001_ VGND VGND VPWR VPWR _00168_ sky130_fd_sc_hd__or2_2
X_09480_ net707 net4272 net659 VGND VGND VPWR VPWR _01233_ sky130_fd_sc_hd__mux2_1
XFILLER_37_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08431_ net1125 _05523_ VGND VGND VPWR VPWR _05524_ sky130_fd_sc_hd__and2_1
XFILLER_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05643_ net30 net1656 VGND VGND VPWR VPWR _03160_ sky130_fd_sc_hd__and2b_1
XFILLER_168_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08362_ net1128 _05477_ VGND VGND VPWR VPWR _05478_ sky130_fd_sc_hd__and2_1
XFILLER_149_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07313_ data_array.data0\[9\]\[52\] net1548 net1452 data_array.data0\[10\]\[52\]
+ VGND VGND VPWR VPWR _04566_ sky130_fd_sc_hd__a22o_1
XFILLER_108_1052 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08293_ net1123 _05431_ VGND VGND VPWR VPWR _05432_ sky130_fd_sc_hd__and2_1
XFILLER_176_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07244_ data_array.data0\[8\]\[46\] net1346 net1252 data_array.data0\[11\]\[46\]
+ _04502_ VGND VGND VPWR VPWR _04503_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_119_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_698 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07175_ net1217 _04435_ _04439_ net1169 VGND VGND VPWR VPWR _04441_ sky130_fd_sc_hd__a22o_1
XFILLER_127_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_882 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06126_ data_array.rdata0\[41\] net1135 net1116 data_array.rdata1\[41\] VGND VGND
+ VPWR VPWR net298 sky130_fd_sc_hd__a22o_1
XFILLER_105_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_184_3920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06057_ net1161 net10 fsm.tag_out1\[11\] net1132 VGND VGND VPWR VPWR _03492_ sky130_fd_sc_hd__a22o_1
XFILLER_133_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_1064 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout334 net335 VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__buf_4
XFILLER_114_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_180_3817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout345 net351 VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__clkbuf_8
XFILLER_86_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout356 net357 VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__buf_4
X_09816_ net945 net3072 net387 VGND VGND VPWR VPWR _01567_ sky130_fd_sc_hd__mux2_1
XFILLER_59_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout367 net368 VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__buf_4
Xfanout378 net379 VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__clkbuf_8
Xfanout389 net393 VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__buf_4
XFILLER_74_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09747_ net700 net3923 net684 VGND VGND VPWR VPWR _01499_ sky130_fd_sc_hd__mux2_1
XFILLER_101_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06959_ data_array.data0\[5\]\[20\] net1603 net1507 data_array.data0\[6\]\[20\] VGND
+ VGND VPWR VPWR _04244_ sky130_fd_sc_hd__a22o_1
XFILLER_100_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09678_ net776 net3294 net605 VGND VGND VPWR VPWR _01430_ sky130_fd_sc_hd__mux2_1
XFILLER_55_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08629_ net706 net4278 net525 VGND VGND VPWR VPWR _00388_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_178_3779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ clknet_leaf_195_clk _00448_ VGND VGND VPWR VPWR tag_array.tag1\[2\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_42_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11571_ clknet_leaf_166_clk _00379_ VGND VGND VPWR VPWR tag_array.tag1\[5\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13310_ clknet_leaf_60_clk _01940_ VGND VGND VPWR VPWR data_array.data0\[10\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_10522_ net857 net4574 net347 VGND VGND VPWR VPWR _02267_ sky130_fd_sc_hd__mux2_1
X_14290_ clknet_leaf_118_clk _02919_ VGND VGND VPWR VPWR data_array.data1\[11\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10453_ net3244 net352 net503 VGND VGND VPWR VPWR _02199_ sky130_fd_sc_hd__mux2_1
X_13241_ clknet_leaf_50_clk _01871_ VGND VGND VPWR VPWR data_array.data0\[11\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_10384_ net1810 net352 net663 VGND VGND VPWR VPWR _02130_ sky130_fd_sc_hd__mux2_1
X_13172_ clknet_leaf_62_clk _00127_ VGND VGND VPWR VPWR data_array.rdata1\[9\] sky130_fd_sc_hd__dfxtp_1
X_12123_ clknet_leaf_146_clk _00931_ VGND VGND VPWR VPWR tag_array.tag0\[12\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_57_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12054_ clknet_leaf_226_clk _00862_ VGND VGND VPWR VPWR data_array.data1\[14\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_123_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11005_ net2019 net982 net336 VGND VGND VPWR VPWR _02749_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout890 _05530_ VGND VGND VPWR VPWR net890 sky130_fd_sc_hd__clkbuf_2
XFILLER_92_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_335 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12956_ clknet_leaf_114_clk _01650_ VGND VGND VPWR VPWR data_array.data0\[13\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_29_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11907_ clknet_leaf_20_clk _00715_ VGND VGND VPWR VPWR data_array.data0\[5\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12887_ clknet_leaf_17_clk _01581_ VGND VGND VPWR VPWR data_array.data0\[12\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
X_11838_ clknet_leaf_127_clk _00646_ VGND VGND VPWR VPWR data_array.data0\[7\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_16_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11769_ clknet_leaf_243_clk _00577_ VGND VGND VPWR VPWR data_array.data0\[8\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_41_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_40_clk clknet_5_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_40_clk sky130_fd_sc_hd__clkbuf_8
X_13508_ clknet_leaf_198_clk _02137_ VGND VGND VPWR VPWR data_array.data1\[0\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_14488_ clknet_leaf_161_clk _03111_ VGND VGND VPWR VPWR tag_array.dirty0\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_158_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload203 clknet_leaf_110_clk VGND VGND VPWR VPWR clkload203/Y sky130_fd_sc_hd__bufinv_16
Xclkload214 clknet_leaf_121_clk VGND VGND VPWR VPWR clkload214/Y sky130_fd_sc_hd__clkinv_4
X_13439_ clknet_leaf_41_clk _02069_ VGND VGND VPWR VPWR data_array.data1\[8\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload225 clknet_leaf_148_clk VGND VGND VPWR VPWR clkload225/Y sky130_fd_sc_hd__inv_6
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload236 clknet_leaf_143_clk VGND VGND VPWR VPWR clkload236/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_161_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08980_ net2026 net1106 net418 VGND VGND VPWR VPWR _00735_ sky130_fd_sc_hd__mux2_1
XFILLER_69_811 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07931_ data_array.data1\[5\]\[44\] net1589 net1493 data_array.data1\[6\]\[44\] VGND
+ VGND VPWR VPWR _05128_ sky130_fd_sc_hd__a22o_1
Xhold2706 data_array.data0\[5\]\[33\] VGND VGND VPWR VPWR net4357 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_138_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2717 data_array.data1\[2\]\[33\] VGND VGND VPWR VPWR net4368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2728 data_array.data0\[11\]\[50\] VGND VGND VPWR VPWR net4379 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_68_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2739 data_array.data1\[10\]\[31\] VGND VGND VPWR VPWR net4390 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07862_ data_array.data1\[0\]\[38\] net1397 net1303 data_array.data1\[3\]\[38\] _05064_
+ VGND VGND VPWR VPWR _05065_ sky130_fd_sc_hd__a221o_1
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09601_ net945 net3109 net394 VGND VGND VPWR VPWR _01353_ sky130_fd_sc_hd__mux2_1
X_06813_ _04110_ _04111_ VGND VGND VPWR VPWR _00060_ sky130_fd_sc_hd__or2_1
X_07793_ data_array.data1\[13\]\[32\] net1521 net1425 data_array.data1\[14\]\[32\]
+ VGND VGND VPWR VPWR _05002_ sky130_fd_sc_hd__a22o_1
XFILLER_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09532_ net698 net4405 net622 VGND VGND VPWR VPWR _01285_ sky130_fd_sc_hd__mux2_1
X_06744_ data_array.data0\[4\]\[0\] net1365 net1271 data_array.data0\[7\]\[0\] _04048_
+ VGND VGND VPWR VPWR _04049_ sky130_fd_sc_hd__a221o_1
XFILLER_3_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09463_ net774 net2829 net653 VGND VGND VPWR VPWR _01216_ sky130_fd_sc_hd__mux2_1
X_06675_ tag_array.tag1\[13\]\[19\] net1579 net1483 tag_array.tag1\[14\]\[19\] VGND
+ VGND VPWR VPWR _03986_ sky130_fd_sc_hd__a22o_1
XFILLER_145_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08414_ net1881 net926 net686 VGND VGND VPWR VPWR _00267_ sky130_fd_sc_hd__mux2_1
XFILLER_12_608 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_05626_ net1649 net1158 VGND VGND VPWR VPWR _03147_ sky130_fd_sc_hd__nand2_2
X_09394_ net1090 net2152 net582 VGND VGND VPWR VPWR _01147_ sky130_fd_sc_hd__mux2_1
X_08345_ net1905 net1018 net688 VGND VGND VPWR VPWR _00244_ sky130_fd_sc_hd__mux2_1
XFILLER_51_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_31_clk clknet_5_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_173_3676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08276_ net3053 net1108 net690 VGND VGND VPWR VPWR _00221_ sky130_fd_sc_hd__mux2_1
XFILLER_164_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_134_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07227_ data_array.data0\[5\]\[44\] net1586 net1490 data_array.data0\[6\]\[44\] VGND
+ VGND VPWR VPWR _04488_ sky130_fd_sc_hd__a22o_1
XFILLER_146_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07158_ data_array.data0\[0\]\[38\] net1396 net1302 data_array.data0\[3\]\[38\] _04424_
+ VGND VGND VPWR VPWR _04425_ sky130_fd_sc_hd__a221o_1
XFILLER_133_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06109_ data_array.rdata0\[24\] net1139 net1115 data_array.rdata1\[24\] VGND VGND
+ VPWR VPWR net279 sky130_fd_sc_hd__a22o_1
XFILLER_65_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07089_ data_array.data0\[13\]\[32\] net1523 net1427 data_array.data0\[14\]\[32\]
+ VGND VGND VPWR VPWR _04362_ sky130_fd_sc_hd__a22o_1
Xfanout1107 _05422_ VGND VGND VPWR VPWR net1107 sky130_fd_sc_hd__buf_1
Xfanout1118 net1119 VGND VGND VPWR VPWR net1118 sky130_fd_sc_hd__clkbuf_4
Xfanout1129 net1130 VGND VGND VPWR VPWR net1129 sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_98_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_98_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_35_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12810_ clknet_leaf_191_clk _01504_ VGND VGND VPWR VPWR tag_array.tag1\[0\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_13790_ clknet_leaf_24_clk _02419_ VGND VGND VPWR VPWR data_array.data1\[2\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_12741_ clknet_leaf_160_clk _01435_ VGND VGND VPWR VPWR tag_array.tag0\[5\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12672_ clknet_leaf_220_clk _01366_ VGND VGND VPWR VPWR data_array.data0\[15\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
X_14411_ clknet_leaf_210_clk _03034_ VGND VGND VPWR VPWR data_array.data1\[10\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11623_ clknet_leaf_168_clk _00431_ VGND VGND VPWR VPWR tag_array.tag1\[3\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_13_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_22_clk clknet_5_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_8
X_14342_ clknet_leaf_121_clk _02971_ VGND VGND VPWR VPWR data_array.data1\[11\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11554_ clknet_leaf_234_clk _00362_ VGND VGND VPWR VPWR tag_array.tag1\[6\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10505_ net926 net2881 net344 VGND VGND VPWR VPWR _02250_ sky130_fd_sc_hd__mux2_1
X_14273_ clknet_leaf_239_clk _02902_ VGND VGND VPWR VPWR data_array.data1\[12\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
X_11485_ clknet_leaf_152_clk _00294_ VGND VGND VPWR VPWR tag_array.valid0\[10\] sky130_fd_sc_hd__dfxtp_1
X_13224_ clknet_leaf_201_clk _00121_ VGND VGND VPWR VPWR data_array.rdata1\[61\] sky130_fd_sc_hd__dfxtp_1
X_10436_ net2061 net908 net662 VGND VGND VPWR VPWR _02182_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13155_ clknet_leaf_140_clk _01849_ VGND VGND VPWR VPWR tag_array.tag1\[8\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_55_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10367_ net733 net4399 net538 VGND VGND VPWR VPWR _02114_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_29_Left_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12106_ clknet_leaf_208_clk _00914_ VGND VGND VPWR VPWR data_array.data1\[14\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10298_ net1961 net969 net633 VGND VGND VPWR VPWR _02045_ sky130_fd_sc_hd__mux2_1
X_13086_ clknet_leaf_216_clk _01780_ VGND VGND VPWR VPWR data_array.data1\[13\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_97_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_89_clk clknet_5_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_89_clk sky130_fd_sc_hd__clkbuf_8
Xfanout1630 net1632 VGND VGND VPWR VPWR net1630 sky130_fd_sc_hd__buf_4
X_12037_ clknet_leaf_90_clk _00845_ VGND VGND VPWR VPWR data_array.data0\[6\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout1641 net1642 VGND VGND VPWR VPWR net1641 sky130_fd_sc_hd__clkbuf_8
XFILLER_38_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13988_ clknet_leaf_30_clk _02617_ VGND VGND VPWR VPWR data_array.data1\[5\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12939_ clknet_leaf_47_clk _01633_ VGND VGND VPWR VPWR data_array.data0\[13\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_38_Left_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06460_ net1221 _03785_ _03789_ net1172 VGND VGND VPWR VPWR _03791_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_138_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_155_3340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06391_ tag_array.tag0\[5\]\[18\] net1597 net1501 tag_array.tag0\[6\]\[18\] VGND
+ VGND VPWR VPWR _03728_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_155_3351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_13_clk clknet_5_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_8
X_08130_ data_array.data1\[0\]\[62\] net1416 net1322 data_array.data1\[3\]\[62\] _05308_
+ VGND VGND VPWR VPWR _05309_ sky130_fd_sc_hd__a221o_1
XFILLER_147_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08061_ data_array.data1\[9\]\[56\] net1532 net1436 data_array.data1\[10\]\[56\]
+ VGND VGND VPWR VPWR _05246_ sky130_fd_sc_hd__a22o_1
XFILLER_105_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07012_ data_array.data0\[13\]\[25\] net1523 net1427 data_array.data0\[14\]\[25\]
+ VGND VGND VPWR VPWR _04292_ sky130_fd_sc_hd__a22o_1
XFILLER_175_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_47_Left_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08963_ net912 net1966 net430 VGND VGND VPWR VPWR _00719_ sky130_fd_sc_hd__mux2_1
Xhold2503 data_array.data1\[9\]\[25\] VGND VGND VPWR VPWR net4154 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2514 data_array.data1\[10\]\[59\] VGND VGND VPWR VPWR net4165 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2525 tag_array.dirty0\[3\] VGND VGND VPWR VPWR net4176 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07914_ data_array.data1\[9\]\[43\] net1568 net1472 data_array.data1\[10\]\[43\]
+ VGND VGND VPWR VPWR _05112_ sky130_fd_sc_hd__a22o_1
Xhold2536 data_array.data0\[11\]\[59\] VGND VGND VPWR VPWR net4187 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1802 data_array.data1\[7\]\[10\] VGND VGND VPWR VPWR net3453 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2547 data_array.data0\[6\]\[25\] VGND VGND VPWR VPWR net4198 sky130_fd_sc_hd__dlygate4sd3_1
X_08894_ net928 net3316 net435 VGND VGND VPWR VPWR _00651_ sky130_fd_sc_hd__mux2_1
Xhold1813 tag_array.tag0\[14\]\[10\] VGND VGND VPWR VPWR net3464 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2558 data_array.data1\[14\]\[5\] VGND VGND VPWR VPWR net4209 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2569 data_array.data0\[11\]\[58\] VGND VGND VPWR VPWR net4220 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1824 tag_array.tag1\[12\]\[3\] VGND VGND VPWR VPWR net3475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1835 tag_array.tag1\[4\]\[23\] VGND VGND VPWR VPWR net3486 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07845_ net1635 _05043_ _05047_ net1209 VGND VGND VPWR VPWR _05050_ sky130_fd_sc_hd__a22o_1
Xhold1846 data_array.data1\[13\]\[56\] VGND VGND VPWR VPWR net3497 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1857 data_array.data1\[11\]\[0\] VGND VGND VPWR VPWR net3508 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1868 data_array.data0\[9\]\[53\] VGND VGND VPWR VPWR net3519 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1879 data_array.data0\[14\]\[13\] VGND VGND VPWR VPWR net3530 sky130_fd_sc_hd__dlygate4sd3_1
X_07776_ data_array.data1\[12\]\[30\] net1394 net1300 data_array.data1\[15\]\[30\]
+ _04986_ VGND VGND VPWR VPWR _04987_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_56_Left_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09515_ net768 net4370 net621 VGND VGND VPWR VPWR _01268_ sky130_fd_sc_hd__mux2_1
XFILLER_37_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06727_ tag_array.tag1\[12\]\[24\] net1372 net1278 tag_array.tag1\[15\]\[24\] _04032_
+ VGND VGND VPWR VPWR _04033_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_175_3716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_175_3727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09446_ net882 net3897 net581 VGND VGND VPWR VPWR _01199_ sky130_fd_sc_hd__mux2_1
X_06658_ net1184 _03965_ _03969_ net1232 VGND VGND VPWR VPWR _03971_ sky130_fd_sc_hd__a22o_1
XFILLER_33_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09377_ net894 net3098 net404 VGND VGND VPWR VPWR _01130_ sky130_fd_sc_hd__mux2_1
XFILLER_149_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06589_ tag_array.tag1\[1\]\[11\] net1575 net1479 tag_array.tag1\[2\]\[11\] VGND
+ VGND VPWR VPWR _03908_ sky130_fd_sc_hd__a22o_1
XFILLER_32_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08328_ net108 net43 net1640 VGND VGND VPWR VPWR _05455_ sky130_fd_sc_hd__mux2_1
XFILLER_149_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08259_ net706 net2573 net805 VGND VGND VPWR VPWR _00217_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_65_Left_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11270_ net951 net3157 net683 VGND VGND VPWR VPWR _03013_ sky130_fd_sc_hd__mux2_1
XFILLER_4_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10221_ net920 net3982 net358 VGND VGND VPWR VPWR _01968_ sky130_fd_sc_hd__mux2_1
XFILLER_161_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10152_ net938 net3614 net366 VGND VGND VPWR VPWR _01900_ sky130_fd_sc_hd__mux2_1
XFILLER_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput290 net290 VGND VGND VPWR VPWR mem_wdata[34] sky130_fd_sc_hd__buf_2
XFILLER_95_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10083_ net1846 net792 net639 VGND VGND VPWR VPWR _01832_ sky130_fd_sc_hd__mux2_1
XFILLER_181_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13911_ clknet_leaf_66_clk _02540_ VGND VGND VPWR VPWR data_array.data1\[4\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_50_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13842_ clknet_leaf_116_clk _02471_ VGND VGND VPWR VPWR data_array.data1\[3\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13773_ clknet_leaf_198_clk _02402_ VGND VGND VPWR VPWR data_array.data1\[2\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10985_ net2388 net1060 net343 VGND VGND VPWR VPWR _02729_ sky130_fd_sc_hd__mux2_1
XFILLER_16_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_861 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12724_ clknet_leaf_109_clk _01418_ VGND VGND VPWR VPWR tag_array.tag0\[7\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12655_ clknet_leaf_218_clk _01349_ VGND VGND VPWR VPWR data_array.data0\[15\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11606_ clknet_leaf_194_clk _00414_ VGND VGND VPWR VPWR tag_array.tag1\[4\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12586_ clknet_leaf_185_clk _01280_ VGND VGND VPWR VPWR tag_array.tag0\[10\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_96_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14325_ clknet_leaf_27_clk _02954_ VGND VGND VPWR VPWR data_array.data1\[11\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
X_11537_ clknet_leaf_191_clk _00345_ VGND VGND VPWR VPWR tag_array.tag1\[6\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_129_679 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold409 data_array.data1\[2\]\[3\] VGND VGND VPWR VPWR net2060 sky130_fd_sc_hd__dlygate4sd3_1
X_14256_ clknet_leaf_122_clk _02885_ VGND VGND VPWR VPWR data_array.data1\[12\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_109_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11468_ clknet_leaf_236_clk _00278_ VGND VGND VPWR VPWR data_array.data0\[0\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_74_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13207_ clknet_leaf_81_clk _00102_ VGND VGND VPWR VPWR data_array.rdata1\[44\] sky130_fd_sc_hd__dfxtp_1
X_10419_ net2947 net978 net668 VGND VGND VPWR VPWR _02165_ sky130_fd_sc_hd__mux2_1
X_14187_ clknet_leaf_244_clk _02816_ VGND VGND VPWR VPWR data_array.data0\[2\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11399_ clknet_leaf_133_clk _00209_ VGND VGND VPWR VPWR tag_array.tag1\[7\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_13138_ clknet_leaf_95_clk _01832_ VGND VGND VPWR VPWR tag_array.tag1\[8\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_112_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13069_ clknet_leaf_122_clk _01763_ VGND VGND VPWR VPWR data_array.data1\[13\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_05960_ data_array.rdata0\[43\] net1658 net1148 VGND VGND VPWR VPWR _03434_ sky130_fd_sc_hd__o21a_1
XFILLER_24_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_2_clk clknet_5_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_8
Xhold1109 tag_array.tag0\[15\]\[2\] VGND VGND VPWR VPWR net2760 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout1460 net1461 VGND VGND VPWR VPWR net1460 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_119_Right_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05891_ data_array.rdata0\[20\] net852 net1149 VGND VGND VPWR VPWR _03388_ sky130_fd_sc_hd__o21a_1
Xfanout1471 net1473 VGND VGND VPWR VPWR net1471 sky130_fd_sc_hd__clkbuf_4
Xfanout1482 net1483 VGND VGND VPWR VPWR net1482 sky130_fd_sc_hd__clkbuf_2
Xfanout1493 net1494 VGND VGND VPWR VPWR net1493 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_109_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07630_ data_array.data1\[1\]\[17\] net1526 net1430 data_array.data1\[2\]\[17\] VGND
+ VGND VPWR VPWR _04854_ sky130_fd_sc_hd__a22o_1
XFILLER_65_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07561_ _04790_ _04791_ VGND VGND VPWR VPWR _00065_ sky130_fd_sc_hd__or2_1
XFILLER_65_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09300_ net778 net3475 net545 VGND VGND VPWR VPWR _01054_ sky130_fd_sc_hd__mux2_1
X_06512_ tag_array.tag1\[5\]\[4\] net1552 net1456 tag_array.tag1\[6\]\[4\] VGND VGND
+ VPWR VPWR _03838_ sky130_fd_sc_hd__a22o_1
X_07492_ data_array.data1\[0\]\[4\] net1393 net1299 data_array.data1\[3\]\[4\] _04728_
+ VGND VGND VPWR VPWR _04729_ sky130_fd_sc_hd__a221o_1
XFILLER_167_708 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09231_ net755 net2392 net646 VGND VGND VPWR VPWR _00985_ sky130_fd_sc_hd__mux2_1
XFILLER_181_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06443_ tag_array.tag0\[0\]\[23\] net1412 net1318 tag_array.tag0\[3\]\[23\] _03774_
+ VGND VGND VPWR VPWR _03775_ sky130_fd_sc_hd__a221o_1
XFILLER_148_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_3624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09162_ net893 net4397 net567 VGND VGND VPWR VPWR _00916_ sky130_fd_sc_hd__mux2_1
X_06374_ tag_array.tag0\[13\]\[17\] net1596 net1500 tag_array.tag0\[14\]\[17\] VGND
+ VGND VPWR VPWR _03712_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_170_3635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08113_ data_array.data1\[12\]\[61\] net1359 net1265 data_array.data1\[15\]\[61\]
+ _05292_ VGND VGND VPWR VPWR _05293_ sky130_fd_sc_hd__a221o_1
X_09093_ net912 net2655 net414 VGND VGND VPWR VPWR _00847_ sky130_fd_sc_hd__mux2_1
XFILLER_119_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08044_ net1218 _05225_ _05229_ net1170 VGND VGND VPWR VPWR _05231_ sky130_fd_sc_hd__a22o_1
XFILLER_119_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_638 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold910 tag_array.tag0\[13\]\[16\] VGND VGND VPWR VPWR net2561 sky130_fd_sc_hd__dlygate4sd3_1
Xhold921 data_array.data0\[4\]\[42\] VGND VGND VPWR VPWR net2572 sky130_fd_sc_hd__dlygate4sd3_1
Xhold932 data_array.data0\[13\]\[3\] VGND VGND VPWR VPWR net2583 sky130_fd_sc_hd__dlygate4sd3_1
Xhold943 data_array.data0\[10\]\[40\] VGND VGND VPWR VPWR net2594 sky130_fd_sc_hd__dlygate4sd3_1
Xhold954 data_array.data1\[4\]\[41\] VGND VGND VPWR VPWR net2605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold965 data_array.data0\[15\]\[40\] VGND VGND VPWR VPWR net2616 sky130_fd_sc_hd__dlygate4sd3_1
Xhold976 data_array.data1\[13\]\[2\] VGND VGND VPWR VPWR net2627 sky130_fd_sc_hd__dlygate4sd3_1
Xhold987 tag_array.tag0\[8\]\[18\] VGND VGND VPWR VPWR net2638 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_168_3586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold998 tag_array.tag0\[8\]\[13\] VGND VGND VPWR VPWR net2649 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_168_3597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09995_ net1106 net3912 net554 VGND VGND VPWR VPWR _01744_ sky130_fd_sc_hd__mux2_1
Xhold2300 data_array.data0\[14\]\[39\] VGND VGND VPWR VPWR net3951 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2311 lru_array.lru_mem\[1\] VGND VGND VPWR VPWR net3962 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2322 tag_array.tag0\[2\]\[10\] VGND VGND VPWR VPWR net3973 sky130_fd_sc_hd__dlygate4sd3_1
X_08946_ net982 net4483 net426 VGND VGND VPWR VPWR _00702_ sky130_fd_sc_hd__mux2_1
XFILLER_9_1050 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2333 data_array.data0\[14\]\[28\] VGND VGND VPWR VPWR net3984 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2344 tag_array.tag0\[13\]\[17\] VGND VGND VPWR VPWR net3995 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2355 tag_array.tag1\[13\]\[9\] VGND VGND VPWR VPWR net4006 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1610 data_array.data0\[9\]\[3\] VGND VGND VPWR VPWR net3261 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1621 tag_array.tag1\[10\]\[17\] VGND VGND VPWR VPWR net3272 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2366 data_array.data1\[11\]\[34\] VGND VGND VPWR VPWR net4017 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1632 tag_array.tag0\[11\]\[24\] VGND VGND VPWR VPWR net3283 sky130_fd_sc_hd__dlygate4sd3_1
X_08877_ net996 net4447 net435 VGND VGND VPWR VPWR _00634_ sky130_fd_sc_hd__mux2_1
Xhold2377 tag_array.tag0\[5\]\[19\] VGND VGND VPWR VPWR net4028 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1643 tag_array.tag0\[5\]\[4\] VGND VGND VPWR VPWR net3294 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2388 data_array.data1\[6\]\[28\] VGND VGND VPWR VPWR net4039 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2399 data_array.data1\[10\]\[26\] VGND VGND VPWR VPWR net4050 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1654 data_array.data0\[13\]\[7\] VGND VGND VPWR VPWR net3305 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1665 data_array.data0\[7\]\[45\] VGND VGND VPWR VPWR net3316 sky130_fd_sc_hd__dlygate4sd3_1
X_07828_ data_array.data1\[5\]\[35\] net1525 net1429 data_array.data1\[6\]\[35\] VGND
+ VGND VPWR VPWR _05034_ sky130_fd_sc_hd__a22o_1
Xhold1676 tag_array.tag1\[7\]\[6\] VGND VGND VPWR VPWR net3327 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1687 data_array.data1\[10\]\[47\] VGND VGND VPWR VPWR net3338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1698 data_array.data1\[8\]\[51\] VGND VGND VPWR VPWR net3349 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07759_ _04970_ _04971_ VGND VGND VPWR VPWR _00084_ sky130_fd_sc_hd__or2_2
XFILLER_44_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10770_ net892 net4172 net493 VGND VGND VPWR VPWR _02515_ sky130_fd_sc_hd__mux2_1
XFILLER_80_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09429_ net951 net4352 net588 VGND VGND VPWR VPWR _01182_ sky130_fd_sc_hd__mux2_1
XFILLER_40_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12440_ clknet_leaf_207_clk _01134_ VGND VGND VPWR VPWR data_array.data0\[14\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
X_12371_ clknet_leaf_2_clk _00048_ VGND VGND VPWR VPWR data_array.rdata0\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_153_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14110_ clknet_leaf_9_clk _02739_ VGND VGND VPWR VPWR data_array.data0\[1\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_11322_ net1004 net4555 net797 VGND VGND VPWR VPWR _03065_ sky130_fd_sc_hd__mux2_1
XFILLER_176_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14041_ clknet_leaf_254_clk _02670_ VGND VGND VPWR VPWR data_array.data1\[6\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_91_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11253_ net1017 net3456 net677 VGND VGND VPWR VPWR _02996_ sky130_fd_sc_hd__mux2_1
XFILLER_69_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10204_ net989 net2707 net359 VGND VGND VPWR VPWR _01951_ sky130_fd_sc_hd__mux2_1
XFILLER_121_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11184_ net1039 net3933 net650 VGND VGND VPWR VPWR _02927_ sky130_fd_sc_hd__mux2_1
XFILLER_122_855 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10135_ net1007 net4582 net362 VGND VGND VPWR VPWR _01883_ sky130_fd_sc_hd__mux2_1
XFILLER_0_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_931 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10066_ net758 net3480 net600 VGND VGND VPWR VPWR _01815_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_89_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13825_ clknet_leaf_220_clk _02454_ VGND VGND VPWR VPWR data_array.data1\[2\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13756_ clknet_leaf_212_clk _02385_ VGND VGND VPWR VPWR data_array.data1\[1\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
X_10968_ net870 net3438 net535 VGND VGND VPWR VPWR _02713_ sky130_fd_sc_hd__mux2_1
XFILLER_31_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12707_ clknet_leaf_107_clk _01401_ VGND VGND VPWR VPWR tag_array.tag0\[7\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_13687_ clknet_leaf_77_clk _02316_ VGND VGND VPWR VPWR data_array.data1\[15\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
X_10899_ net890 net3470 net515 VGND VGND VPWR VPWR _02644_ sky130_fd_sc_hd__mux2_1
XFILLER_176_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12638_ clknet_leaf_128_clk _01332_ VGND VGND VPWR VPWR data_array.data0\[15\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_100_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12569_ clknet_leaf_164_clk _01263_ VGND VGND VPWR VPWR tag_array.tag0\[10\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_157_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14308_ clknet_leaf_30_clk _02937_ VGND VGND VPWR VPWR data_array.data1\[11\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_06090_ data_array.rdata0\[5\] net1136 net1117 data_array.rdata1\[5\] VGND VGND VPWR
+ VPWR net318 sky130_fd_sc_hd__a22o_1
XFILLER_172_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold206 data_array.data0\[2\]\[26\] VGND VGND VPWR VPWR net1857 sky130_fd_sc_hd__dlygate4sd3_1
Xhold217 data_array.data0\[4\]\[26\] VGND VGND VPWR VPWR net1868 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold228 data_array.data0\[1\]\[31\] VGND VGND VPWR VPWR net1879 sky130_fd_sc_hd__dlygate4sd3_1
X_14239_ clknet_leaf_204_clk _02868_ VGND VGND VPWR VPWR data_array.data1\[12\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold239 tag_array.tag1\[0\]\[15\] VGND VGND VPWR VPWR net1890 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout708 _05407_ VGND VGND VPWR VPWR net708 sky130_fd_sc_hd__clkbuf_2
Xfanout719 net721 VGND VGND VPWR VPWR net719 sky130_fd_sc_hd__clkbuf_2
X_08800_ net2322 net1046 net444 VGND VGND VPWR VPWR _00558_ sky130_fd_sc_hd__mux2_1
X_09780_ net1089 net2394 net388 VGND VGND VPWR VPWR _01531_ sky130_fd_sc_hd__mux2_1
XFILLER_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06992_ data_array.data0\[1\]\[23\] net1556 net1460 data_array.data0\[2\]\[23\] VGND
+ VGND VPWR VPWR _04274_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_146_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08731_ net2719 net700 net476 VGND VGND VPWR VPWR _00490_ sky130_fd_sc_hd__mux2_1
X_05943_ data_array.rdata1\[37\] net830 net839 VGND VGND VPWR VPWR _03423_ sky130_fd_sc_hd__a21o_1
XFILLER_67_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_163_3494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1290 net1291 VGND VGND VPWR VPWR net1290 sky130_fd_sc_hd__clkbuf_4
X_08662_ net775 net4019 net494 VGND VGND VPWR VPWR _00421_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05874_ data_array.rdata1\[14\] net833 net842 VGND VGND VPWR VPWR _03377_ sky130_fd_sc_hd__a21o_1
XFILLER_27_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07613_ data_array.data1\[0\]\[15\] net1394 net1300 data_array.data1\[3\]\[15\] _04838_
+ VGND VGND VPWR VPWR _04839_ sky130_fd_sc_hd__a221o_1
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08593_ net750 net3965 net535 VGND VGND VPWR VPWR _00352_ sky130_fd_sc_hd__mux2_1
XFILLER_41_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07544_ data_array.data1\[13\]\[9\] net1581 net1485 data_array.data1\[14\]\[9\] VGND
+ VGND VPWR VPWR _04776_ sky130_fd_sc_hd__a22o_1
XFILLER_14_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07475_ data_array.data1\[12\]\[3\] net1384 net1290 data_array.data1\[15\]\[3\] _04712_
+ VGND VGND VPWR VPWR _04713_ sky130_fd_sc_hd__a221o_1
X_09214_ net722 net3995 net631 VGND VGND VPWR VPWR _00968_ sky130_fd_sc_hd__mux2_1
XFILLER_179_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06426_ net1211 _03753_ _03757_ net1637 VGND VGND VPWR VPWR _03760_ sky130_fd_sc_hd__a22o_1
XFILLER_50_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09145_ net960 net2983 net566 VGND VGND VPWR VPWR _00899_ sky130_fd_sc_hd__mux2_1
XFILLER_182_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06357_ tag_array.tag0\[8\]\[15\] net1402 net1308 tag_array.tag0\[11\]\[15\] _03696_
+ VGND VGND VPWR VPWR _03697_ sky130_fd_sc_hd__a221o_1
XFILLER_136_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09076_ net982 net4560 net410 VGND VGND VPWR VPWR _00830_ sky130_fd_sc_hd__mux2_1
X_06288_ tag_array.tag0\[1\]\[9\] net1598 net1502 tag_array.tag0\[2\]\[9\] VGND VGND
+ VPWR VPWR _03634_ sky130_fd_sc_hd__a22o_1
XFILLER_162_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08027_ data_array.data1\[0\]\[53\] net1333 net1239 data_array.data1\[3\]\[53\] _05214_
+ VGND VGND VPWR VPWR _05215_ sky130_fd_sc_hd__a221o_1
Xhold740 data_array.data1\[8\]\[4\] VGND VGND VPWR VPWR net2391 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold751 data_array.data0\[4\]\[45\] VGND VGND VPWR VPWR net2402 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold762 data_array.data1\[8\]\[33\] VGND VGND VPWR VPWR net2413 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold773 data_array.data0\[0\]\[25\] VGND VGND VPWR VPWR net2424 sky130_fd_sc_hd__dlygate4sd3_1
Xhold784 data_array.data0\[4\]\[33\] VGND VGND VPWR VPWR net2435 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_118_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold795 tag_array.tag0\[11\]\[16\] VGND VGND VPWR VPWR net2446 sky130_fd_sc_hd__dlygate4sd3_1
X_09978_ net916 net2994 net376 VGND VGND VPWR VPWR _01727_ sky130_fd_sc_hd__mux2_1
Xhold2130 data_array.data0\[3\]\[16\] VGND VGND VPWR VPWR net3781 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2141 tag_array.tag0\[7\]\[8\] VGND VGND VPWR VPWR net3792 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_46 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2152 data_array.data0\[9\]\[40\] VGND VGND VPWR VPWR net3803 sky130_fd_sc_hd__dlygate4sd3_1
X_08929_ net1048 net2286 net430 VGND VGND VPWR VPWR _00685_ sky130_fd_sc_hd__mux2_1
Xhold2163 data_array.data0\[3\]\[50\] VGND VGND VPWR VPWR net3814 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2174 tag_array.tag0\[7\]\[6\] VGND VGND VPWR VPWR net3825 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2185 data_array.data1\[7\]\[20\] VGND VGND VPWR VPWR net3836 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1440 data_array.data0\[14\]\[33\] VGND VGND VPWR VPWR net3091 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1451 lru_array.lru_mem\[14\] VGND VGND VPWR VPWR net3102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2196 data_array.data1\[14\]\[20\] VGND VGND VPWR VPWR net3847 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11940_ clknet_leaf_50_clk _00748_ VGND VGND VPWR VPWR data_array.data0\[4\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_55_22 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1462 tag_array.tag0\[14\]\[8\] VGND VGND VPWR VPWR net3113 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1473 data_array.data1\[9\]\[20\] VGND VGND VPWR VPWR net3124 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1484 tag_array.tag1\[6\]\[0\] VGND VGND VPWR VPWR net3135 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1495 data_array.data0\[8\]\[54\] VGND VGND VPWR VPWR net3146 sky130_fd_sc_hd__dlygate4sd3_1
X_11871_ clknet_leaf_62_clk _00679_ VGND VGND VPWR VPWR data_array.data0\[5\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_73_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13610_ clknet_leaf_243_clk _02239_ VGND VGND VPWR VPWR data_array.data0\[9\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
X_10822_ net1960 net942 net509 VGND VGND VPWR VPWR _02567_ sky130_fd_sc_hd__mux2_1
XFILLER_38_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13541_ clknet_leaf_74_clk _02170_ VGND VGND VPWR VPWR data_array.data1\[0\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1055 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10753_ net963 net4132 net493 VGND VGND VPWR VPWR _02498_ sky130_fd_sc_hd__mux2_1
XFILLER_40_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13472_ clknet_leaf_179_clk _02102_ VGND VGND VPWR VPWR tag_array.tag0\[15\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_10684_ net3888 net980 net478 VGND VGND VPWR VPWR _02429_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12423_ clknet_leaf_260_clk _01117_ VGND VGND VPWR VPWR data_array.data0\[14\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_154_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12354_ clknet_leaf_118_clk _00029_ VGND VGND VPWR VPWR data_array.rdata0\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11305_ net1075 net4434 net801 VGND VGND VPWR VPWR _03048_ sky130_fd_sc_hd__mux2_1
X_12285_ clknet_leaf_141_clk _01043_ VGND VGND VPWR VPWR tag_array.tag1\[13\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14024_ clknet_leaf_227_clk _02653_ VGND VGND VPWR VPWR data_array.data1\[6\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_11236_ net1087 net3111 net673 VGND VGND VPWR VPWR _02979_ sky130_fd_sc_hd__mux2_1
XFILLER_106_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11167_ net1107 net3844 net648 VGND VGND VPWR VPWR _02910_ sky130_fd_sc_hd__mux2_1
XFILLER_121_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10118_ net1073 net3690 net367 VGND VGND VPWR VPWR _01866_ sky130_fd_sc_hd__mux2_1
X_11098_ net1909 net868 net335 VGND VGND VPWR VPWR _02841_ sky130_fd_sc_hd__mux2_1
XFILLER_110_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10049_ net891 net3036 net556 VGND VGND VPWR VPWR _01798_ sky130_fd_sc_hd__mux2_1
XFILLER_48_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_141_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13808_ clknet_leaf_123_clk _02437_ VGND VGND VPWR VPWR data_array.data1\[2\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_102_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_11_Left_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13739_ clknet_leaf_257_clk _02368_ VGND VGND VPWR VPWR data_array.data1\[1\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07260_ data_array.data0\[1\]\[47\] net1577 net1481 data_array.data0\[2\]\[47\] VGND
+ VGND VPWR VPWR _04518_ sky130_fd_sc_hd__a22o_1
X_06211_ tag_array.tag0\[5\]\[2\] net1560 net1464 tag_array.tag0\[6\]\[2\] VGND VGND
+ VPWR VPWR _03564_ sky130_fd_sc_hd__a22o_1
X_07191_ data_array.data0\[4\]\[41\] net1337 net1243 data_array.data0\[7\]\[41\] _04454_
+ VGND VGND VPWR VPWR _04455_ sky130_fd_sc_hd__a221o_1
XFILLER_117_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06142_ data_array.rdata0\[57\] net1136 net1117 data_array.rdata1\[57\] VGND VGND
+ VPWR VPWR net315 sky130_fd_sc_hd__a22o_1
X_06073_ net1161 net19 fsm.tag_out1\[19\] net1133 VGND VGND VPWR VPWR _03500_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_148_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09901_ net866 net3017 net381 VGND VGND VPWR VPWR _01651_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_6_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_3534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout505 net506 VGND VGND VPWR VPWR net505 sky130_fd_sc_hd__buf_4
XFILLER_113_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout516 net517 VGND VGND VPWR VPWR net516 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_6_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09832_ net881 net3683 net389 VGND VGND VPWR VPWR _01583_ sky130_fd_sc_hd__mux2_1
Xfanout527 net530 VGND VGND VPWR VPWR net527 sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_171_Right_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout538 net540 VGND VGND VPWR VPWR net538 sky130_fd_sc_hd__buf_4
Xfanout549 net553 VGND VGND VPWR VPWR net549 sky130_fd_sc_hd__buf_4
XFILLER_101_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09763_ net2767 net735 net665 VGND VGND VPWR VPWR _01515_ sky130_fd_sc_hd__mux2_1
XFILLER_112_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06975_ data_array.data0\[4\]\[21\] net1365 net1271 data_array.data0\[7\]\[21\] _04258_
+ VGND VGND VPWR VPWR _04259_ sky130_fd_sc_hd__a221o_1
X_08714_ net2015 net766 net469 VGND VGND VPWR VPWR _00473_ sky130_fd_sc_hd__mux2_1
XFILLER_39_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05926_ net123 net1156 _03411_ _03410_ VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__a22o_1
X_09694_ net712 net3288 net605 VGND VGND VPWR VPWR _01446_ sky130_fd_sc_hd__mux2_1
XFILLER_27_636 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08645_ net3405 net743 net511 VGND VGND VPWR VPWR _00404_ sky130_fd_sc_hd__mux2_1
X_05857_ net161 net1151 _03364_ _03365_ VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__a22o_1
XFILLER_81_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08576_ net812 _05587_ VGND VGND VPWR VPWR _05603_ sky130_fd_sc_hd__and2_1
XFILLER_109_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05788_ _03136_ fsm.tag_out1\[2\] _03277_ VGND VGND VPWR VPWR _03305_ sky130_fd_sc_hd__a21o_1
X_07527_ net1227 _04755_ _04759_ net1179 VGND VGND VPWR VPWR _04761_ sky130_fd_sc_hd__a22o_1
XFILLER_148_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_875 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07458_ data_array.data1\[5\]\[1\] net1520 net1424 data_array.data1\[6\]\[1\] VGND
+ VGND VPWR VPWR _04698_ sky130_fd_sc_hd__a22o_1
XFILLER_168_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06409_ tag_array.tag0\[5\]\[20\] net1558 net1462 tag_array.tag0\[6\]\[20\] VGND
+ VGND VPWR VPWR _03744_ sky130_fd_sc_hd__a22o_1
XFILLER_183_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07389_ data_array.data0\[0\]\[59\] net1379 net1285 data_array.data0\[3\]\[59\] _04634_
+ VGND VGND VPWR VPWR _04635_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_40_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09128_ net1031 net3847 net576 VGND VGND VPWR VPWR _00882_ sky130_fd_sc_hd__mux2_1
XFILLER_157_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09059_ net1048 net2518 net414 VGND VGND VPWR VPWR _00813_ sky130_fd_sc_hd__mux2_1
XFILLER_155_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_724 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12070_ clknet_leaf_218_clk _00878_ VGND VGND VPWR VPWR data_array.data1\[14\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold570 lru_array.lru_mem\[6\] VGND VGND VPWR VPWR net2221 sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 data_array.data0\[8\]\[27\] VGND VGND VPWR VPWR net2232 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold592 tag_array.tag1\[14\]\[18\] VGND VGND VPWR VPWR net2243 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_663 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11021_ net2219 net916 net342 VGND VGND VPWR VPWR _02765_ sky130_fd_sc_hd__mux2_1
XFILLER_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12972_ clknet_leaf_155_clk _01666_ VGND VGND VPWR VPWR tag_array.tag0\[4\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_46_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1270 data_array.data1\[8\]\[18\] VGND VGND VPWR VPWR net2921 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11923_ clknet_leaf_207_clk _00731_ VGND VGND VPWR VPWR data_array.data0\[5\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1281 tag_array.tag0\[14\]\[1\] VGND VGND VPWR VPWR net2932 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1292 data_array.data1\[6\]\[6\] VGND VGND VPWR VPWR net2943 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11854_ clknet_leaf_12_clk _00662_ VGND VGND VPWR VPWR data_array.data0\[7\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_64_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_680 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10805_ net2633 net1008 net502 VGND VGND VPWR VPWR _02550_ sky130_fd_sc_hd__mux2_1
X_11785_ clknet_leaf_3_clk _00593_ VGND VGND VPWR VPWR data_array.data0\[8\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
X_13524_ clknet_leaf_228_clk _02153_ VGND VGND VPWR VPWR data_array.data1\[0\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_10736_ net1030 net2896 net500 VGND VGND VPWR VPWR _02481_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13455_ clknet_leaf_165_clk _02085_ VGND VGND VPWR VPWR tag_array.tag0\[1\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_10667_ net1743 net1051 net484 VGND VGND VPWR VPWR _02412_ sky130_fd_sc_hd__mux2_1
XFILLER_127_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12406_ clknet_leaf_34_clk _01100_ VGND VGND VPWR VPWR data_array.data0\[14\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_13386_ clknet_leaf_268_clk _02016_ VGND VGND VPWR VPWR data_array.data1\[8\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10598_ net1872 net1070 net475 VGND VGND VPWR VPWR _02343_ sky130_fd_sc_hd__mux2_1
XFILLER_154_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12337_ clknet_leaf_67_clk _00010_ VGND VGND VPWR VPWR data_array.rdata0\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_56_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12268_ clknet_leaf_96_clk _01026_ VGND VGND VPWR VPWR tag_array.tag1\[13\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_123_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14007_ clknet_leaf_78_clk _02636_ VGND VGND VPWR VPWR data_array.data1\[5\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
X_11219_ net899 net4586 net648 VGND VGND VPWR VPWR _02962_ sky130_fd_sc_hd__mux2_1
XFILLER_123_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12199_ clknet_leaf_183_clk _00152_ VGND VGND VPWR VPWR fsm.tag_out0\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_143_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06760_ data_array.data0\[12\]\[2\] net1338 net1244 data_array.data0\[15\]\[2\] _04062_
+ VGND VGND VPWR VPWR _04063_ sky130_fd_sc_hd__a221o_1
XFILLER_110_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05711_ _03182_ _03184_ _03200_ fsm.valid0 VGND VGND VPWR VPWR _03228_ sky130_fd_sc_hd__or4b_1
X_06691_ net1222 _03995_ _03999_ net1173 VGND VGND VPWR VPWR _04001_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_121_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08430_ net146 net81 net1643 VGND VGND VPWR VPWR _05523_ sky130_fd_sc_hd__mux2_1
X_05642_ _03155_ _03156_ _03157_ _03158_ VGND VGND VPWR VPWR _03159_ sky130_fd_sc_hd__or4_1
XFILLER_52_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08361_ net120 net55 net1640 VGND VGND VPWR VPWR _05477_ sky130_fd_sc_hd__mux2_1
XFILLER_108_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07312_ data_array.data0\[4\]\[52\] net1355 net1261 data_array.data0\[7\]\[52\] _04564_
+ VGND VGND VPWR VPWR _04565_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_22_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08292_ net159 net94 net1638 VGND VGND VPWR VPWR _05431_ sky130_fd_sc_hd__mux2_1
XFILLER_20_845 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07243_ data_array.data0\[9\]\[46\] net1537 net1441 data_array.data0\[10\]\[46\]
+ VGND VGND VPWR VPWR _04502_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_119_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07174_ net1619 _04433_ _04437_ net1193 VGND VGND VPWR VPWR _04440_ sky130_fd_sc_hd__a22o_1
XFILLER_11_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_266_clk clknet_5_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_266_clk
+ sky130_fd_sc_hd__clkbuf_8
X_06125_ data_array.rdata0\[40\] _03477_ net1119 data_array.rdata1\[40\] VGND VGND
+ VPWR VPWR net297 sky130_fd_sc_hd__a22o_1
XFILLER_133_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_184_3910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_184_3921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06056_ fsm.tag_out0\[10\] net1121 _03491_ VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_132_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_180_3818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout335 _03133_ VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__buf_4
XFILLER_99_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_1076 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout346 net347 VGND VGND VPWR VPWR net346 sky130_fd_sc_hd__buf_4
X_09815_ net949 net2954 net392 VGND VGND VPWR VPWR _01566_ sky130_fd_sc_hd__mux2_1
Xfanout357 net361 VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__clkbuf_4
XFILLER_87_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout368 net369 VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__clkbuf_8
Xfanout379 net385 VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__buf_4
XFILLER_87_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09746_ net702 net2115 net678 VGND VGND VPWR VPWR _01498_ sky130_fd_sc_hd__mux2_1
X_06958_ data_array.data0\[12\]\[20\] net1419 net1325 data_array.data0\[15\]\[20\]
+ _04242_ VGND VGND VPWR VPWR _04243_ sky130_fd_sc_hd__a221o_1
XFILLER_39_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05909_ data_array.rdata0\[26\] net846 net1142 VGND VGND VPWR VPWR _03400_ sky130_fd_sc_hd__o21a_1
XFILLER_55_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09677_ net779 net3169 net605 VGND VGND VPWR VPWR _01429_ sky130_fd_sc_hd__mux2_1
XFILLER_36_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06889_ net1219 _04175_ _04179_ net1171 VGND VGND VPWR VPWR _04181_ sky130_fd_sc_hd__a22o_1
XFILLER_28_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08628_ net710 net4360 net515 VGND VGND VPWR VPWR _00387_ sky130_fd_sc_hd__mux2_1
X_08559_ net719 net2672 net584 VGND VGND VPWR VPWR _00327_ sky130_fd_sc_hd__mux2_1
XFILLER_35_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11570_ clknet_leaf_33_clk _00378_ VGND VGND VPWR VPWR tag_array.tag1\[5\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10521_ net861 net3237 net351 VGND VGND VPWR VPWR _02266_ sky130_fd_sc_hd__mux2_1
XFILLER_161_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13240_ clknet_leaf_192_clk _01870_ VGND VGND VPWR VPWR data_array.data0\[11\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_10452_ net352 net4556 net519 VGND VGND VPWR VPWR _02198_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_257_clk clknet_5_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_257_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13171_ clknet_leaf_15_clk _00126_ VGND VGND VPWR VPWR data_array.rdata1\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_124_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10383_ net352 net4282 net675 VGND VGND VPWR VPWR _02129_ sky130_fd_sc_hd__mux2_1
XFILLER_163_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12122_ clknet_leaf_181_clk _00930_ VGND VGND VPWR VPWR tag_array.tag0\[12\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12053_ clknet_leaf_226_clk _00861_ VGND VGND VPWR VPWR data_array.data0\[6\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_77_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11004_ net1879 net986 net342 VGND VGND VPWR VPWR _02748_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout880 net881 VGND VGND VPWR VPWR net880 sky130_fd_sc_hd__clkbuf_2
Xfanout891 _05530_ VGND VGND VPWR VPWR net891 sky130_fd_sc_hd__buf_1
XFILLER_46_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12955_ clknet_leaf_51_clk _01649_ VGND VGND VPWR VPWR data_array.data0\[13\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_29_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11906_ clknet_leaf_87_clk _00714_ VGND VGND VPWR VPWR data_array.data0\[5\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_179_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12886_ clknet_leaf_219_clk _01580_ VGND VGND VPWR VPWR data_array.data0\[12\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_45_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11837_ clknet_leaf_235_clk _00645_ VGND VGND VPWR VPWR data_array.data0\[7\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_159_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11768_ clknet_leaf_10_clk _00576_ VGND VGND VPWR VPWR data_array.data0\[8\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
X_13507_ clknet_leaf_69_clk _02136_ VGND VGND VPWR VPWR data_array.data1\[0\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10719_ net1098 net3915 net496 VGND VGND VPWR VPWR _02464_ sky130_fd_sc_hd__mux2_1
XFILLER_146_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14487_ clknet_leaf_161_clk _03110_ VGND VGND VPWR VPWR tag_array.dirty0\[6\] sky130_fd_sc_hd__dfxtp_1
X_11699_ clknet_leaf_100_clk _00507_ VGND VGND VPWR VPWR tag_array.tag1\[15\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_173_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload204 clknet_leaf_111_clk VGND VGND VPWR VPWR clkload204/Y sky130_fd_sc_hd__clkinv_2
Xclkload215 clknet_leaf_122_clk VGND VGND VPWR VPWR clkload215/X sky130_fd_sc_hd__clkbuf_4
X_13438_ clknet_leaf_202_clk _02068_ VGND VGND VPWR VPWR data_array.data1\[8\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
Xrebuffer1 _03194_ VGND VGND VPWR VPWR net1652 sky130_fd_sc_hd__dlygate4sd1_1
Xclkload226 clknet_leaf_150_clk VGND VGND VPWR VPWR clkload226/Y sky130_fd_sc_hd__inv_12
Xclkload237 clknet_leaf_133_clk VGND VGND VPWR VPWR clkload237/Y sky130_fd_sc_hd__inv_6
Xclkbuf_leaf_248_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_248_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_155_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13369_ clknet_leaf_231_clk _01999_ VGND VGND VPWR VPWR tag_array.tag0\[2\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_77_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07930_ data_array.data1\[12\]\[44\] net1398 net1304 data_array.data1\[15\]\[44\]
+ _05126_ VGND VGND VPWR VPWR _05127_ sky130_fd_sc_hd__a221o_1
XFILLER_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2707 data_array.data1\[7\]\[29\] VGND VGND VPWR VPWR net4358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2718 tag_array.tag0\[6\]\[4\] VGND VGND VPWR VPWR net4369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2729 tag_array.tag0\[4\]\[20\] VGND VGND VPWR VPWR net4380 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07861_ data_array.data1\[1\]\[38\] net1588 net1492 data_array.data1\[2\]\[38\] VGND
+ VGND VPWR VPWR _05064_ sky130_fd_sc_hd__a22o_1
X_09600_ net949 net2616 net400 VGND VGND VPWR VPWR _01352_ sky130_fd_sc_hd__mux2_1
X_06812_ net1213 _04105_ _04109_ net1165 VGND VGND VPWR VPWR _04111_ sky130_fd_sc_hd__a22o_1
X_07792_ _05000_ _05001_ VGND VGND VPWR VPWR _00088_ sky130_fd_sc_hd__or2_1
X_09531_ net705 net2961 net621 VGND VGND VPWR VPWR _01284_ sky130_fd_sc_hd__mux2_1
XFILLER_3_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06743_ data_array.data0\[5\]\[0\] net1555 net1459 data_array.data0\[6\]\[0\] VGND
+ VGND VPWR VPWR _04048_ sky130_fd_sc_hd__a22o_1
XFILLER_83_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09462_ net778 net3645 net653 VGND VGND VPWR VPWR _01215_ sky130_fd_sc_hd__mux2_1
XFILLER_92_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06674_ tag_array.tag1\[4\]\[19\] net1386 net1292 tag_array.tag1\[7\]\[19\] _03984_
+ VGND VGND VPWR VPWR _03985_ sky130_fd_sc_hd__a221o_1
X_08413_ net1123 _05511_ VGND VGND VPWR VPWR _05512_ sky130_fd_sc_hd__and2_1
X_05625_ net1649 net1160 VGND VGND VPWR VPWR _03146_ sky130_fd_sc_hd__and2_1
XFILLER_184_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09393_ net1095 net3709 net586 VGND VGND VPWR VPWR _01146_ sky130_fd_sc_hd__mux2_1
X_08344_ net1126 _05465_ VGND VGND VPWR VPWR _05466_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_173_3677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08275_ net1130 _05419_ VGND VGND VPWR VPWR _05420_ sky130_fd_sc_hd__and2_1
X_07226_ data_array.data0\[12\]\[44\] net1395 net1301 data_array.data0\[15\]\[44\]
+ _04486_ VGND VGND VPWR VPWR _04487_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_134_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_239_clk clknet_5_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_239_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_121_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07157_ data_array.data0\[1\]\[38\] net1585 net1489 data_array.data0\[2\]\[38\] VGND
+ VGND VPWR VPWR _04424_ sky130_fd_sc_hd__a22o_1
X_06108_ data_array.rdata0\[23\] net1137 net1118 data_array.rdata1\[23\] VGND VGND
+ VPWR VPWR net278 sky130_fd_sc_hd__a22o_1
X_07088_ _04360_ _04361_ VGND VGND VPWR VPWR _00024_ sky130_fd_sc_hd__or2_2
XFILLER_161_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06039_ net1159 net32 fsm.tag_out1\[2\] net1131 VGND VGND VPWR VPWR _03483_ sky130_fd_sc_hd__a22o_1
XFILLER_133_588 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1108 _05420_ VGND VGND VPWR VPWR net1108 sky130_fd_sc_hd__clkbuf_2
XFILLER_114_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1119 _03480_ VGND VGND VPWR VPWR net1119 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_35_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09729_ net772 net2416 net683 VGND VGND VPWR VPWR _01481_ sky130_fd_sc_hd__mux2_1
XFILLER_16_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12740_ clknet_leaf_144_clk _01434_ VGND VGND VPWR VPWR tag_array.tag0\[5\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12671_ clknet_leaf_3_clk _01365_ VGND VGND VPWR VPWR data_array.data0\[15\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_179_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14410_ clknet_leaf_120_clk _03033_ VGND VGND VPWR VPWR data_array.data1\[10\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11622_ clknet_leaf_134_clk _00430_ VGND VGND VPWR VPWR tag_array.tag1\[3\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14341_ clknet_leaf_210_clk _02970_ VGND VGND VPWR VPWR data_array.data1\[11\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
X_11553_ clknet_leaf_98_clk _00361_ VGND VGND VPWR VPWR tag_array.tag1\[6\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10504_ net929 net3393 net345 VGND VGND VPWR VPWR _02249_ sky130_fd_sc_hd__mux2_1
XFILLER_128_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14272_ clknet_leaf_21_clk _02901_ VGND VGND VPWR VPWR data_array.data1\[12\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
X_11484_ clknet_leaf_151_clk _00293_ VGND VGND VPWR VPWR tag_array.valid0\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_59_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13223_ clknet_leaf_119_clk _00120_ VGND VGND VPWR VPWR data_array.rdata1\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_171_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10435_ net1962 net914 net668 VGND VGND VPWR VPWR _02181_ sky130_fd_sc_hd__mux2_1
XFILLER_137_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13154_ clknet_leaf_136_clk _01848_ VGND VGND VPWR VPWR tag_array.tag1\[8\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_10366_ net737 net2857 net538 VGND VGND VPWR VPWR _02113_ sky130_fd_sc_hd__mux2_1
XFILLER_88_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12105_ clknet_leaf_4_clk _00913_ VGND VGND VPWR VPWR data_array.data1\[14\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13085_ clknet_leaf_82_clk _01779_ VGND VGND VPWR VPWR data_array.data1\[13\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10297_ net1971 net974 net633 VGND VGND VPWR VPWR _02044_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12036_ clknet_leaf_244_clk _00844_ VGND VGND VPWR VPWR data_array.data0\[6\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout1620 net1627 VGND VGND VPWR VPWR net1620 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_72_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1631 net1632 VGND VGND VPWR VPWR net1631 sky130_fd_sc_hd__buf_4
Xfanout1642 net98 VGND VGND VPWR VPWR net1642 sky130_fd_sc_hd__buf_8
XFILLER_93_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13987_ clknet_leaf_219_clk _02616_ VGND VGND VPWR VPWR data_array.data1\[5\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_46_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12938_ clknet_leaf_93_clk _01632_ VGND VGND VPWR VPWR data_array.data0\[13\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_138_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12869_ clknet_leaf_219_clk _01563_ VGND VGND VPWR VPWR data_array.data0\[12\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_138_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06390_ tag_array.tag0\[8\]\[18\] net1374 net1280 tag_array.tag0\[11\]\[18\] _03726_
+ VGND VGND VPWR VPWR _03727_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_155_3341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_3352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08060_ data_array.data1\[4\]\[56\] net1340 net1246 data_array.data1\[7\]\[56\] _05244_
+ VGND VGND VPWR VPWR _05245_ sky130_fd_sc_hd__a221o_1
XFILLER_175_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07011_ _04290_ _04291_ VGND VGND VPWR VPWR _00016_ sky130_fd_sc_hd__or2_1
XFILLER_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08962_ net917 net2952 net430 VGND VGND VPWR VPWR _00718_ sky130_fd_sc_hd__mux2_1
XFILLER_102_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2504 data_array.data0\[5\]\[38\] VGND VGND VPWR VPWR net4155 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2515 data_array.data1\[5\]\[38\] VGND VGND VPWR VPWR net4166 sky130_fd_sc_hd__dlygate4sd3_1
X_07913_ _05110_ _05111_ VGND VGND VPWR VPWR _00100_ sky130_fd_sc_hd__or2_1
Xhold2526 data_array.data0\[6\]\[22\] VGND VGND VPWR VPWR net4177 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_124_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2537 data_array.data1\[14\]\[29\] VGND VGND VPWR VPWR net4188 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08893_ net932 net3756 net440 VGND VGND VPWR VPWR _00650_ sky130_fd_sc_hd__mux2_1
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1803 data_array.data0\[14\]\[8\] VGND VGND VPWR VPWR net3454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2548 data_array.data0\[14\]\[18\] VGND VGND VPWR VPWR net4199 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1814 data_array.data1\[9\]\[39\] VGND VGND VPWR VPWR net3465 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2559 tag_array.tag1\[7\]\[11\] VGND VGND VPWR VPWR net4210 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1825 data_array.data1\[7\]\[14\] VGND VGND VPWR VPWR net3476 sky130_fd_sc_hd__dlygate4sd3_1
X_07844_ data_array.data1\[0\]\[36\] net1414 net1320 data_array.data1\[3\]\[36\] _05048_
+ VGND VGND VPWR VPWR _05049_ sky130_fd_sc_hd__a221o_1
XFILLER_151_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1836 tag_array.tag0\[9\]\[2\] VGND VGND VPWR VPWR net3487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1847 data_array.data0\[12\]\[43\] VGND VGND VPWR VPWR net3498 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1858 data_array.data1\[14\]\[35\] VGND VGND VPWR VPWR net3509 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1869 data_array.data1\[5\]\[18\] VGND VGND VPWR VPWR net3520 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07775_ data_array.data1\[13\]\[30\] net1583 net1487 data_array.data1\[14\]\[30\]
+ VGND VGND VPWR VPWR _04986_ sky130_fd_sc_hd__a22o_1
Xclone6 net835 VGND VGND VPWR VPWR net1657 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_3_Left_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09514_ net771 net2758 net623 VGND VGND VPWR VPWR _01267_ sky130_fd_sc_hd__mux2_1
X_06726_ tag_array.tag1\[13\]\[24\] net1562 net1466 tag_array.tag1\[14\]\[24\] VGND
+ VGND VPWR VPWR _04032_ sky130_fd_sc_hd__a22o_1
XFILLER_24_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_175_3717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_175_3728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09445_ net887 net3473 net580 VGND VGND VPWR VPWR _01198_ sky130_fd_sc_hd__mux2_1
X_06657_ net1210 _03963_ _03967_ net1636 VGND VGND VPWR VPWR _03970_ sky130_fd_sc_hd__a22o_1
XFILLER_52_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09376_ net896 net4463 net402 VGND VGND VPWR VPWR _01129_ sky130_fd_sc_hd__mux2_1
X_06588_ tag_array.tag1\[12\]\[11\] net1385 net1291 tag_array.tag1\[15\]\[11\] _03906_
+ VGND VGND VPWR VPWR _03907_ sky130_fd_sc_hd__a221o_1
XFILLER_21_940 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08327_ net1729 net1042 net689 VGND VGND VPWR VPWR _00238_ sky130_fd_sc_hd__mux2_1
X_08258_ fsm.tag_out1\[21\] net818 net810 fsm.tag_out0\[21\] _05406_ VGND VGND VPWR
+ VPWR _05407_ sky130_fd_sc_hd__a221o_2
XFILLER_165_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_494 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07209_ _04470_ _04471_ VGND VGND VPWR VPWR _00036_ sky130_fd_sc_hd__or2_1
X_08189_ net1644 net831 _05358_ VGND VGND VPWR VPWR _05359_ sky130_fd_sc_hd__and3_1
XFILLER_152_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10220_ net926 net3044 net354 VGND VGND VPWR VPWR _01967_ sky130_fd_sc_hd__mux2_1
XFILLER_165_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_363 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10151_ net940 net2714 net368 VGND VGND VPWR VPWR _01899_ sky130_fd_sc_hd__mux2_1
Xoutput280 net280 VGND VGND VPWR VPWR mem_wdata[25] sky130_fd_sc_hd__buf_2
XFILLER_160_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput291 net291 VGND VGND VPWR VPWR mem_wdata[35] sky130_fd_sc_hd__buf_2
X_10082_ net694 net2702 net601 VGND VGND VPWR VPWR _01831_ sky130_fd_sc_hd__mux2_1
XFILLER_88_962 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13910_ clknet_leaf_42_clk _02539_ VGND VGND VPWR VPWR data_array.data1\[4\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_101_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13841_ clknet_leaf_60_clk _02470_ VGND VGND VPWR VPWR data_array.data1\[3\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13772_ clknet_leaf_69_clk _02401_ VGND VGND VPWR VPWR data_array.data1\[2\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_10984_ net1973 net1064 net342 VGND VGND VPWR VPWR _02728_ sky130_fd_sc_hd__mux2_1
XFILLER_55_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12723_ clknet_leaf_157_clk _01417_ VGND VGND VPWR VPWR tag_array.tag0\[7\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_71_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12654_ clknet_leaf_114_clk _01348_ VGND VGND VPWR VPWR data_array.data0\[15\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
X_11605_ clknet_leaf_100_clk _00413_ VGND VGND VPWR VPWR tag_array.tag1\[4\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_96_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12585_ clknet_leaf_108_clk _01279_ VGND VGND VPWR VPWR tag_array.tag0\[10\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_96_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14324_ clknet_leaf_80_clk _02953_ VGND VGND VPWR VPWR data_array.data1\[11\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
X_11536_ clknet_leaf_31_clk _00344_ VGND VGND VPWR VPWR tag_array.tag1\[6\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_117_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_80 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14255_ clknet_leaf_240_clk _02884_ VGND VGND VPWR VPWR data_array.data1\[12\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
X_11467_ clknet_leaf_12_clk _00277_ VGND VGND VPWR VPWR data_array.data0\[0\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_74_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1051 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13206_ clknet_leaf_49_clk _00101_ VGND VGND VPWR VPWR data_array.rdata1\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_143_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10418_ net2177 net980 net661 VGND VGND VPWR VPWR _02164_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14186_ clknet_leaf_11_clk _02815_ VGND VGND VPWR VPWR data_array.data0\[2\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
X_11398_ clknet_leaf_166_clk _00208_ VGND VGND VPWR VPWR tag_array.tag1\[7\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_180_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13137_ clknet_leaf_190_clk _01831_ VGND VGND VPWR VPWR tag_array.tag0\[3\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_10349_ net705 net4459 net594 VGND VGND VPWR VPWR _02096_ sky130_fd_sc_hd__mux2_1
XFILLER_140_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13068_ clknet_leaf_67_clk _01762_ VGND VGND VPWR VPWR data_array.data1\[13\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_97_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1450 net1458 VGND VGND VPWR VPWR net1450 sky130_fd_sc_hd__buf_2
X_12019_ clknet_leaf_52_clk _00827_ VGND VGND VPWR VPWR data_array.data0\[6\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout1461 net1470 VGND VGND VPWR VPWR net1461 sky130_fd_sc_hd__clkbuf_2
X_05890_ net109 net1155 _03386_ _03387_ VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__a22o_1
XFILLER_66_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1472 net1473 VGND VGND VPWR VPWR net1472 sky130_fd_sc_hd__clkbuf_4
XFILLER_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1483 net1495 VGND VGND VPWR VPWR net1483 sky130_fd_sc_hd__clkbuf_4
Xfanout1494 net1495 VGND VGND VPWR VPWR net1494 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_109_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07560_ net1183 _04785_ _04789_ net1233 VGND VGND VPWR VPWR _04791_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06511_ tag_array.tag1\[12\]\[4\] net1362 net1268 tag_array.tag1\[15\]\[4\] _03836_
+ VGND VGND VPWR VPWR _03837_ sky130_fd_sc_hd__a221o_1
XFILLER_80_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07491_ data_array.data1\[1\]\[4\] net1583 net1487 data_array.data1\[2\]\[4\] VGND
+ VGND VPWR VPWR _04728_ sky130_fd_sc_hd__a22o_1
XFILLER_94_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09230_ net759 net3113 net647 VGND VGND VPWR VPWR _00984_ sky130_fd_sc_hd__mux2_1
X_06442_ tag_array.tag0\[1\]\[23\] net1602 net1506 tag_array.tag0\[2\]\[23\] VGND
+ VGND VPWR VPWR _03774_ sky130_fd_sc_hd__a22o_1
XFILLER_166_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09161_ net898 net4570 net566 VGND VGND VPWR VPWR _00915_ sky130_fd_sc_hd__mux2_1
X_06373_ _03710_ _03711_ VGND VGND VPWR VPWR _00138_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_170_3625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08112_ data_array.data1\[13\]\[61\] net1550 net1454 data_array.data1\[14\]\[61\]
+ VGND VGND VPWR VPWR _05292_ sky130_fd_sc_hd__a22o_1
XFILLER_148_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09092_ net917 net3851 net415 VGND VGND VPWR VPWR _00846_ sky130_fd_sc_hd__mux2_1
XFILLER_119_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08043_ net1621 _05223_ _05227_ net1195 VGND VGND VPWR VPWR _05230_ sky130_fd_sc_hd__a22o_1
XFILLER_162_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold900 data_array.data0\[5\]\[26\] VGND VGND VPWR VPWR net2551 sky130_fd_sc_hd__dlygate4sd3_1
Xhold911 data_array.data0\[7\]\[20\] VGND VGND VPWR VPWR net2562 sky130_fd_sc_hd__dlygate4sd3_1
Xhold922 tag_array.tag1\[7\]\[21\] VGND VGND VPWR VPWR net2573 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold933 tag_array.tag0\[6\]\[12\] VGND VGND VPWR VPWR net2584 sky130_fd_sc_hd__dlygate4sd3_1
Xhold944 data_array.data1\[3\]\[15\] VGND VGND VPWR VPWR net2595 sky130_fd_sc_hd__dlygate4sd3_1
Xhold955 data_array.data0\[1\]\[0\] VGND VGND VPWR VPWR net2606 sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 tag_array.tag1\[14\]\[4\] VGND VGND VPWR VPWR net2617 sky130_fd_sc_hd__dlygate4sd3_1
Xhold977 data_array.data1\[1\]\[54\] VGND VGND VPWR VPWR net2628 sky130_fd_sc_hd__dlygate4sd3_1
Xhold988 data_array.data0\[7\]\[60\] VGND VGND VPWR VPWR net2639 sky130_fd_sc_hd__dlygate4sd3_1
X_09994_ net1111 net3746 net559 VGND VGND VPWR VPWR _01743_ sky130_fd_sc_hd__mux2_1
XFILLER_142_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_168_3587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold999 data_array.data0\[13\]\[37\] VGND VGND VPWR VPWR net2650 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_168_3598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2301 data_array.data0\[14\]\[12\] VGND VGND VPWR VPWR net3952 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2312 data_array.data0\[15\]\[13\] VGND VGND VPWR VPWR net3963 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08945_ net987 net4533 net433 VGND VGND VPWR VPWR _00701_ sky130_fd_sc_hd__mux2_1
Xhold2323 tag_array.tag0\[5\]\[15\] VGND VGND VPWR VPWR net3974 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2334 tag_array.tag1\[0\]\[23\] VGND VGND VPWR VPWR net3985 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1600 tag_array.tag0\[0\]\[1\] VGND VGND VPWR VPWR net3251 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2345 tag_array.tag0\[4\]\[3\] VGND VGND VPWR VPWR net3996 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1611 data_array.data0\[12\]\[18\] VGND VGND VPWR VPWR net3262 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2356 tag_array.tag0\[9\]\[17\] VGND VGND VPWR VPWR net4007 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1622 data_array.data1\[7\]\[47\] VGND VGND VPWR VPWR net3273 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2367 data_array.data1\[12\]\[16\] VGND VGND VPWR VPWR net4018 sky130_fd_sc_hd__dlygate4sd3_1
X_08876_ net1003 net4351 net436 VGND VGND VPWR VPWR _00633_ sky130_fd_sc_hd__mux2_1
XFILLER_151_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2378 data_array.data0\[12\]\[1\] VGND VGND VPWR VPWR net4029 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1633 data_array.data1\[10\]\[52\] VGND VGND VPWR VPWR net3284 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1644 data_array.data1\[9\]\[44\] VGND VGND VPWR VPWR net3295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2389 data_array.data1\[13\]\[11\] VGND VGND VPWR VPWR net4040 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1655 data_array.data1\[9\]\[32\] VGND VGND VPWR VPWR net3306 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07827_ data_array.data1\[12\]\[35\] net1335 net1241 data_array.data1\[15\]\[35\]
+ _05032_ VGND VGND VPWR VPWR _05033_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_4_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1666 data_array.data1\[15\]\[38\] VGND VGND VPWR VPWR net3317 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1677 data_array.data0\[6\]\[4\] VGND VGND VPWR VPWR net3328 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1688 data_array.data0\[12\]\[37\] VGND VGND VPWR VPWR net3339 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_71_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1699 tag_array.tag1\[13\]\[11\] VGND VGND VPWR VPWR net3350 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07758_ net1175 _04965_ _04969_ net1223 VGND VGND VPWR VPWR _04971_ sky130_fd_sc_hd__a22o_1
XFILLER_37_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06709_ tag_array.tag1\[8\]\[22\] net1360 net1266 tag_array.tag1\[11\]\[22\] _04016_
+ VGND VGND VPWR VPWR _04017_ sky130_fd_sc_hd__a221o_1
X_07689_ data_array.data1\[5\]\[22\] net1533 net1437 data_array.data1\[6\]\[22\] VGND
+ VGND VPWR VPWR _04908_ sky130_fd_sc_hd__a22o_1
X_09428_ net952 net3465 net581 VGND VGND VPWR VPWR _01181_ sky130_fd_sc_hd__mux2_1
XFILLER_100_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09359_ net964 net3727 net408 VGND VGND VPWR VPWR _01112_ sky130_fd_sc_hd__mux2_1
XFILLER_60_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12370_ clknet_leaf_212_clk _00047_ VGND VGND VPWR VPWR data_array.rdata0\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_165_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_16__f_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_5_16__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_11321_ net1008 net4474 net795 VGND VGND VPWR VPWR _03064_ sky130_fd_sc_hd__mux2_1
XFILLER_153_414 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14040_ clknet_leaf_214_clk _02669_ VGND VGND VPWR VPWR data_array.data1\[6\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_91_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11252_ net1021 net4538 net675 VGND VGND VPWR VPWR _02995_ sky130_fd_sc_hd__mux2_1
XFILLER_4_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10203_ net992 net4329 net359 VGND VGND VPWR VPWR _01950_ sky130_fd_sc_hd__mux2_1
XFILLER_69_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11183_ net1040 net3857 net649 VGND VGND VPWR VPWR _02926_ sky130_fd_sc_hd__mux2_1
XFILLER_106_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10134_ net1009 net4219 net362 VGND VGND VPWR VPWR _01882_ sky130_fd_sc_hd__mux2_1
XFILLER_122_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10065_ net763 net3891 net601 VGND VGND VPWR VPWR _01814_ sky130_fd_sc_hd__mux2_1
XFILLER_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2890 data_array.data0\[10\]\[63\] VGND VGND VPWR VPWR net4541 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_36_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13824_ clknet_leaf_9_clk _02453_ VGND VGND VPWR VPWR data_array.data1\[2\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_391 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13755_ clknet_leaf_4_clk _02384_ VGND VGND VPWR VPWR data_array.data1\[1\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_67_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10967_ net875 net4486 net531 VGND VGND VPWR VPWR _02712_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12706_ clknet_leaf_185_clk _01400_ VGND VGND VPWR VPWR tag_array.tag0\[8\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_10898_ net892 net2985 net516 VGND VGND VPWR VPWR _02643_ sky130_fd_sc_hd__mux2_1
X_13686_ clknet_leaf_6_clk _02315_ VGND VGND VPWR VPWR data_array.data1\[15\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12637_ clknet_leaf_59_clk _01331_ VGND VGND VPWR VPWR data_array.data0\[15\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_169_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12568_ clknet_leaf_106_clk _01262_ VGND VGND VPWR VPWR tag_array.tag0\[10\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_152_Right_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14307_ clknet_leaf_221_clk _02936_ VGND VGND VPWR VPWR data_array.data1\[11\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_11519_ clknet_leaf_187_clk _00327_ VGND VGND VPWR VPWR tag_array.tag1\[9\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_12499_ clknet_leaf_5_clk _01193_ VGND VGND VPWR VPWR data_array.data1\[9\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold207 data_array.data1\[0\]\[57\] VGND VGND VPWR VPWR net1858 sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 data_array.data1\[8\]\[62\] VGND VGND VPWR VPWR net1869 sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 tag_array.tag1\[8\]\[6\] VGND VGND VPWR VPWR net1880 sky130_fd_sc_hd__dlygate4sd3_1
X_14238_ clknet_leaf_241_clk _02867_ VGND VGND VPWR VPWR data_array.data1\[12\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_14169_ clknet_leaf_249_clk _02798_ VGND VGND VPWR VPWR data_array.data0\[2\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout709 _05407_ VGND VGND VPWR VPWR net709 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_84_Left_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06991_ data_array.data0\[12\]\[23\] net1371 net1277 data_array.data0\[15\]\[23\]
+ _04272_ VGND VGND VPWR VPWR _04273_ sky130_fd_sc_hd__a221o_1
XFILLER_112_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08730_ net2196 net702 net469 VGND VGND VPWR VPWR _00489_ sky130_fd_sc_hd__mux2_1
X_05942_ data_array.rdata0\[37\] net848 net1144 VGND VGND VPWR VPWR _03422_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_163_3495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1280 net1281 VGND VGND VPWR VPWR net1280 sky130_fd_sc_hd__clkbuf_4
X_08661_ net778 net4163 net494 VGND VGND VPWR VPWR _00420_ sky130_fd_sc_hd__mux2_1
Xfanout1291 net1294 VGND VGND VPWR VPWR net1291 sky130_fd_sc_hd__clkbuf_4
XFILLER_22_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05873_ data_array.rdata0\[14\] net851 net1148 VGND VGND VPWR VPWR _03376_ sky130_fd_sc_hd__o21a_1
XFILLER_38_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07612_ data_array.data1\[1\]\[15\] net1584 net1488 data_array.data1\[2\]\[15\] VGND
+ VGND VPWR VPWR _04838_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_124_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08592_ net756 net4567 net535 VGND VGND VPWR VPWR _00351_ sky130_fd_sc_hd__mux2_1
X_07543_ data_array.data1\[4\]\[9\] net1389 net1295 data_array.data1\[7\]\[9\] _04774_
+ VGND VGND VPWR VPWR _04775_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_93_Left_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07474_ data_array.data1\[13\]\[3\] net1574 net1478 data_array.data1\[14\]\[3\] VGND
+ VGND VPWR VPWR _04712_ sky130_fd_sc_hd__a22o_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09213_ net727 net2561 net631 VGND VGND VPWR VPWR _00967_ sky130_fd_sc_hd__mux2_1
X_06425_ tag_array.tag0\[0\]\[21\] net1407 net1313 tag_array.tag0\[3\]\[21\] _03758_
+ VGND VGND VPWR VPWR _03759_ sky130_fd_sc_hd__a221o_1
XFILLER_22_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09144_ net967 net2800 net574 VGND VGND VPWR VPWR _00898_ sky130_fd_sc_hd__mux2_1
X_06356_ tag_array.tag0\[9\]\[15\] net1594 net1498 tag_array.tag0\[10\]\[15\] VGND
+ VGND VPWR VPWR _03696_ sky130_fd_sc_hd__a22o_1
XFILLER_148_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09075_ net986 net4564 net416 VGND VGND VPWR VPWR _00829_ sky130_fd_sc_hd__mux2_1
XFILLER_147_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06287_ tag_array.tag0\[12\]\[9\] net1409 net1315 tag_array.tag0\[15\]\[9\] _03632_
+ VGND VGND VPWR VPWR _03633_ sky130_fd_sc_hd__a221o_1
X_08026_ data_array.data1\[1\]\[53\] net1524 net1428 data_array.data1\[2\]\[53\] VGND
+ VGND VPWR VPWR _05214_ sky130_fd_sc_hd__a22o_1
Xhold730 data_array.data0\[0\]\[16\] VGND VGND VPWR VPWR net2381 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold741 tag_array.tag0\[14\]\[9\] VGND VGND VPWR VPWR net2392 sky130_fd_sc_hd__dlygate4sd3_1
Xhold752 data_array.data1\[2\]\[57\] VGND VGND VPWR VPWR net2403 sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 lru_array.lru_mem\[9\] VGND VGND VPWR VPWR net2414 sky130_fd_sc_hd__dlygate4sd3_1
Xhold774 data_array.data0\[9\]\[61\] VGND VGND VPWR VPWR net2425 sky130_fd_sc_hd__dlygate4sd3_1
Xhold785 data_array.data0\[1\]\[60\] VGND VGND VPWR VPWR net2436 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_118_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold796 tag_array.tag1\[3\]\[19\] VGND VGND VPWR VPWR net2447 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09977_ net921 net3907 net375 VGND VGND VPWR VPWR _01726_ sky130_fd_sc_hd__mux2_1
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2120 tag_array.tag1\[6\]\[21\] VGND VGND VPWR VPWR net3771 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2131 data_array.data0\[15\]\[51\] VGND VGND VPWR VPWR net3782 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2142 data_array.data1\[6\]\[22\] VGND VGND VPWR VPWR net3793 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_58 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08928_ net1052 net3489 net431 VGND VGND VPWR VPWR _00684_ sky130_fd_sc_hd__mux2_1
Xhold2153 data_array.data1\[7\]\[49\] VGND VGND VPWR VPWR net3804 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2164 data_array.data0\[6\]\[45\] VGND VGND VPWR VPWR net3815 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2175 data_array.data0\[11\]\[22\] VGND VGND VPWR VPWR net3826 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1430 tag_array.tag1\[8\]\[12\] VGND VGND VPWR VPWR net3081 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2186 data_array.data0\[7\]\[4\] VGND VGND VPWR VPWR net3837 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1441 data_array.data0\[6\]\[13\] VGND VGND VPWR VPWR net3092 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1452 data_array.data1\[11\]\[54\] VGND VGND VPWR VPWR net3103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2197 data_array.data0\[15\]\[29\] VGND VGND VPWR VPWR net3848 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1463 data_array.data1\[4\]\[38\] VGND VGND VPWR VPWR net3114 sky130_fd_sc_hd__dlygate4sd3_1
X_08859_ net1068 net2513 net440 VGND VGND VPWR VPWR _00616_ sky130_fd_sc_hd__mux2_1
Xhold1474 data_array.data0\[5\]\[52\] VGND VGND VPWR VPWR net3125 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1485 tag_array.tag0\[14\]\[13\] VGND VGND VPWR VPWR net3136 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1496 tag_array.tag1\[15\]\[3\] VGND VGND VPWR VPWR net3147 sky130_fd_sc_hd__dlygate4sd3_1
X_11870_ clknet_leaf_14_clk _00678_ VGND VGND VPWR VPWR data_array.data0\[5\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_169_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10821_ net2605 net944 net502 VGND VGND VPWR VPWR _02566_ sky130_fd_sc_hd__mux2_1
XFILLER_77_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10752_ net965 net2426 net497 VGND VGND VPWR VPWR _02497_ sky130_fd_sc_hd__mux2_1
X_13540_ clknet_leaf_214_clk _02169_ VGND VGND VPWR VPWR data_array.data1\[0\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_45_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1067 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13471_ clknet_leaf_170_clk _02101_ VGND VGND VPWR VPWR tag_array.tag0\[15\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_41_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10683_ net3501 net984 net483 VGND VGND VPWR VPWR _02428_ sky130_fd_sc_hd__mux2_1
XFILLER_125_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12422_ clknet_leaf_124_clk _01116_ VGND VGND VPWR VPWR data_array.data0\[14\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_71_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12353_ clknet_leaf_256_clk _00028_ VGND VGND VPWR VPWR data_array.rdata0\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_126_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11304_ net1078 net3524 net796 VGND VGND VPWR VPWR _03047_ sky130_fd_sc_hd__mux2_1
X_12284_ clknet_leaf_136_clk _01042_ VGND VGND VPWR VPWR tag_array.tag1\[13\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14023_ clknet_leaf_204_clk _02652_ VGND VGND VPWR VPWR data_array.data1\[5\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11235_ net1091 net2147 net677 VGND VGND VPWR VPWR _02978_ sky130_fd_sc_hd__mux2_1
XFILLER_135_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11166_ net1111 net3508 net654 VGND VGND VPWR VPWR _02909_ sky130_fd_sc_hd__mux2_1
XFILLER_84_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10117_ net1076 net4189 net363 VGND VGND VPWR VPWR _01865_ sky130_fd_sc_hd__mux2_1
XFILLER_110_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11097_ net2444 net872 net334 VGND VGND VPWR VPWR _02840_ sky130_fd_sc_hd__mux2_1
XFILLER_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10048_ net893 net2569 net555 VGND VGND VPWR VPWR _01797_ sky130_fd_sc_hd__mux2_1
XFILLER_48_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_69_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_106_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold90 data_array.data1\[0\]\[10\] VGND VGND VPWR VPWR net1741 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_64_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13807_ clknet_leaf_240_clk _02436_ VGND VGND VPWR VPWR data_array.data1\[2\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11999_ clknet_leaf_62_clk _00807_ VGND VGND VPWR VPWR data_array.data0\[6\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_82_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13738_ clknet_leaf_10_clk _02367_ VGND VGND VPWR VPWR data_array.data1\[1\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_82_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_859 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13669_ clknet_leaf_39_clk _02298_ VGND VGND VPWR VPWR data_array.data1\[15\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_06210_ tag_array.tag0\[8\]\[2\] net1369 net1275 tag_array.tag0\[11\]\[2\] _03562_
+ VGND VGND VPWR VPWR _03563_ sky130_fd_sc_hd__a221o_1
X_07190_ data_array.data0\[5\]\[41\] net1527 net1431 data_array.data0\[6\]\[41\] VGND
+ VGND VPWR VPWR _04454_ sky130_fd_sc_hd__a22o_1
XFILLER_118_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06141_ data_array.rdata0\[56\] net1135 net1112 data_array.rdata1\[56\] VGND VGND
+ VPWR VPWR net314 sky130_fd_sc_hd__a22o_1
XFILLER_129_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06072_ fsm.tag_out0\[18\] _03478_ _03499_ VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__a21o_1
XFILLER_117_469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09900_ net868 net2933 net384 VGND VGND VPWR VPWR _01650_ sky130_fd_sc_hd__mux2_1
XFILLER_116_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_165_3524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout506 net513 VGND VGND VPWR VPWR net506 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_165_3535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout517 net518 VGND VGND VPWR VPWR net517 sky130_fd_sc_hd__clkbuf_8
X_09831_ net885 net3593 net387 VGND VGND VPWR VPWR _01582_ sky130_fd_sc_hd__mux2_1
Xfanout528 net529 VGND VGND VPWR VPWR net528 sky130_fd_sc_hd__buf_4
Xfanout539 net540 VGND VGND VPWR VPWR net539 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_182_3860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09762_ net2135 net741 net672 VGND VGND VPWR VPWR _01514_ sky130_fd_sc_hd__mux2_1
X_06974_ data_array.data0\[5\]\[21\] net1555 net1459 data_array.data0\[6\]\[21\] VGND
+ VGND VPWR VPWR _04258_ sky130_fd_sc_hd__a22o_1
X_08713_ net1812 net772 net475 VGND VGND VPWR VPWR _00472_ sky130_fd_sc_hd__mux2_1
X_05925_ data_array.rdata1\[31\] net833 net842 VGND VGND VPWR VPWR _03411_ sky130_fd_sc_hd__a21o_1
X_09693_ net716 net4028 net606 VGND VGND VPWR VPWR _01445_ sky130_fd_sc_hd__mux2_1
XFILLER_39_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08644_ net2486 net746 net507 VGND VGND VPWR VPWR _00403_ sky130_fd_sc_hd__mux2_1
X_05856_ data_array.rdata1\[8\] net829 net838 VGND VGND VPWR VPWR _03365_ sky130_fd_sc_hd__a21o_1
XFILLER_148_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08575_ net1727 net482 VGND VGND VPWR VPWR _00338_ sky130_fd_sc_hd__or2_1
XFILLER_42_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_05787_ _03136_ fsm.tag_out1\[2\] fsm.valid1 VGND VGND VPWR VPWR _03304_ sky130_fd_sc_hd__o21ai_1
XFILLER_41_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07526_ net1631 _04753_ _04757_ net1205 VGND VGND VPWR VPWR _04760_ sky130_fd_sc_hd__a22o_1
XFILLER_23_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07457_ data_array.data1\[8\]\[1\] net1330 net1236 data_array.data1\[11\]\[1\] _04696_
+ VGND VGND VPWR VPWR _04697_ sky130_fd_sc_hd__a221o_1
X_06408_ tag_array.tag0\[12\]\[20\] net1369 net1276 tag_array.tag0\[15\]\[20\] _03742_
+ VGND VGND VPWR VPWR _03743_ sky130_fd_sc_hd__a221o_1
X_07388_ data_array.data0\[1\]\[59\] net1570 net1474 data_array.data0\[2\]\[59\] VGND
+ VGND VPWR VPWR _04634_ sky130_fd_sc_hd__a22o_1
XFILLER_176_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09127_ net1035 net4031 net574 VGND VGND VPWR VPWR _00881_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06339_ net1232 _03675_ _03679_ net1184 VGND VGND VPWR VPWR _03681_ sky130_fd_sc_hd__a22o_1
XFILLER_136_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09058_ net1052 net4347 net415 VGND VGND VPWR VPWR _00812_ sky130_fd_sc_hd__mux2_1
XFILLER_68_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08009_ data_array.data1\[0\]\[51\] net1332 net1238 data_array.data1\[3\]\[51\] _05198_
+ VGND VGND VPWR VPWR _05199_ sky130_fd_sc_hd__a221o_1
XFILLER_2_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold560 data_array.data0\[4\]\[11\] VGND VGND VPWR VPWR net2211 sky130_fd_sc_hd__dlygate4sd3_1
Xhold571 data_array.data0\[8\]\[3\] VGND VGND VPWR VPWR net2222 sky130_fd_sc_hd__dlygate4sd3_1
Xhold582 tag_array.tag1\[7\]\[18\] VGND VGND VPWR VPWR net2233 sky130_fd_sc_hd__dlygate4sd3_1
X_11020_ net2070 net920 net342 VGND VGND VPWR VPWR _02764_ sky130_fd_sc_hd__mux2_1
XFILLER_173_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold593 data_array.data0\[2\]\[47\] VGND VGND VPWR VPWR net2244 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12971_ clknet_leaf_165_clk _01665_ VGND VGND VPWR VPWR tag_array.tag0\[4\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_85_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1260 data_array.data1\[11\]\[52\] VGND VGND VPWR VPWR net2911 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1271 data_array.data1\[3\]\[51\] VGND VGND VPWR VPWR net2922 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1282 data_array.data0\[13\]\[60\] VGND VGND VPWR VPWR net2933 sky130_fd_sc_hd__dlygate4sd3_1
X_11922_ clknet_leaf_111_clk _00730_ VGND VGND VPWR VPWR data_array.data0\[5\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1293 data_array.data0\[9\]\[52\] VGND VGND VPWR VPWR net2944 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11853_ clknet_leaf_14_clk _00661_ VGND VGND VPWR VPWR data_array.data0\[7\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_64_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10804_ net2148 net1015 net508 VGND VGND VPWR VPWR _02549_ sky130_fd_sc_hd__mux2_1
X_11784_ clknet_leaf_241_clk _00592_ VGND VGND VPWR VPWR data_array.data0\[8\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
X_13523_ clknet_leaf_130_clk _02152_ VGND VGND VPWR VPWR data_array.data1\[0\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_10735_ net1034 net2301 net497 VGND VGND VPWR VPWR _02480_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_24_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10666_ net2980 net1054 net483 VGND VGND VPWR VPWR _02411_ sky130_fd_sc_hd__mux2_1
X_13454_ clknet_leaf_105_clk _02084_ VGND VGND VPWR VPWR tag_array.tag0\[1\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_174_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_149_Left_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12405_ clknet_leaf_176_clk _01099_ VGND VGND VPWR VPWR data_array.data0\[14\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_13385_ clknet_leaf_198_clk _02015_ VGND VGND VPWR VPWR data_array.data1\[8\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10597_ net1730 net1074 net472 VGND VGND VPWR VPWR _02342_ sky130_fd_sc_hd__mux2_1
XFILLER_182_851 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12336_ clknet_leaf_15_clk _00009_ VGND VGND VPWR VPWR data_array.rdata0\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12267_ clknet_leaf_188_clk _01025_ VGND VGND VPWR VPWR tag_array.tag1\[14\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_141_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11218_ net901 net2911 net652 VGND VGND VPWR VPWR _02961_ sky130_fd_sc_hd__mux2_1
X_14006_ clknet_leaf_261_clk _02635_ VGND VGND VPWR VPWR data_array.data1\[5\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_68_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12198_ clknet_leaf_146_clk _00151_ VGND VGND VPWR VPWR fsm.tag_out0\[5\] sky130_fd_sc_hd__dfxtp_2
XFILLER_150_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_143_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11149_ net923 net4276 net550 VGND VGND VPWR VPWR _02892_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_143_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_158_Left_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_160_3432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05710_ _03156_ _03158_ _03203_ VGND VGND VPWR VPWR _03227_ sky130_fd_sc_hd__or3_1
X_06690_ net1625 _03993_ _03997_ net1200 VGND VGND VPWR VPWR _04000_ sky130_fd_sc_hd__a22o_1
XFILLER_64_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05641_ net7 fsm.tag_out0\[8\] VGND VGND VPWR VPWR _03158_ sky130_fd_sc_hd__xor2_1
XFILLER_17_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08360_ net2345 net996 net687 VGND VGND VPWR VPWR _00249_ sky130_fd_sc_hd__mux2_1
X_07311_ data_array.data0\[5\]\[52\] net1545 net1449 data_array.data0\[6\]\[52\] VGND
+ VGND VPWR VPWR _04564_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_22_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_3394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08291_ net1985 net1088 net688 VGND VGND VPWR VPWR _00226_ sky130_fd_sc_hd__mux2_1
XFILLER_32_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_167_Left_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07242_ _04500_ _04501_ VGND VGND VPWR VPWR _00039_ sky130_fd_sc_hd__or2_1
XFILLER_20_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07173_ data_array.data0\[4\]\[39\] net1348 net1254 data_array.data0\[7\]\[39\] _04438_
+ VGND VGND VPWR VPWR _04439_ sky130_fd_sc_hd__a221o_1
XFILLER_157_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06124_ data_array.rdata0\[39\] net1135 net1116 data_array.rdata1\[39\] VGND VGND
+ VPWR VPWR net295 sky130_fd_sc_hd__a22o_1
XFILLER_145_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_184_3900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06055_ net1163 net9 fsm.tag_out1\[10\] net1132 VGND VGND VPWR VPWR _03491_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_184_3911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_184_3922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_180_3819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_176_Left_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout336 net340 VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__buf_4
XFILLER_98_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout347 net351 VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__clkbuf_4
X_09814_ net955 net4121 net389 VGND VGND VPWR VPWR _01565_ sky130_fd_sc_hd__mux2_1
XFILLER_143_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout358 net360 VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__buf_4
Xfanout369 _03128_ VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__clkbuf_8
XFILLER_87_868 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09745_ net707 net3203 net684 VGND VGND VPWR VPWR _01497_ sky130_fd_sc_hd__mux2_1
X_06957_ data_array.data0\[13\]\[20\] net1609 net1513 data_array.data0\[14\]\[20\]
+ VGND VGND VPWR VPWR _04242_ sky130_fd_sc_hd__a22o_1
XFILLER_95_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05908_ net116 net1150 _03398_ _03399_ VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__a22o_1
XFILLER_39_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06888_ net1197 _04173_ _04177_ net1622 VGND VGND VPWR VPWR _04180_ sky130_fd_sc_hd__a22o_1
X_09676_ net784 net3759 net605 VGND VGND VPWR VPWR _01428_ sky130_fd_sc_hd__mux2_1
XFILLER_28_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05839_ net121 net1151 _03352_ _03353_ VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__a22o_1
X_08627_ net714 net3448 net522 VGND VGND VPWR VPWR _00386_ sky130_fd_sc_hd__mux2_1
XFILLER_160_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08558_ net725 net4105 net588 VGND VGND VPWR VPWR _00326_ sky130_fd_sc_hd__mux2_1
XFILLER_51_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07509_ data_array.data1\[1\]\[6\] net1519 net1423 data_array.data1\[2\]\[6\] VGND
+ VGND VPWR VPWR _04744_ sky130_fd_sc_hd__a22o_1
XFILLER_167_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08489_ net824 net813 net855 _05561_ VGND VGND VPWR VPWR _05563_ sky130_fd_sc_hd__or4b_1
XFILLER_168_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10520_ net867 net2425 net346 VGND VGND VPWR VPWR _02265_ sky130_fd_sc_hd__mux2_1
XFILLER_161_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10451_ net352 net4381 net531 VGND VGND VPWR VPWR _02197_ sky130_fd_sc_hd__mux2_1
X_13170_ clknet_leaf_81_clk _00125_ VGND VGND VPWR VPWR data_array.rdata1\[7\] sky130_fd_sc_hd__dfxtp_1
X_10382_ net352 net3477 net650 VGND VGND VPWR VPWR _02128_ sky130_fd_sc_hd__mux2_1
X_12121_ clknet_leaf_179_clk _00929_ VGND VGND VPWR VPWR tag_array.tag0\[12\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12052_ clknet_leaf_109_clk _00860_ VGND VGND VPWR VPWR data_array.data0\[6\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold390 data_array.data1\[8\]\[53\] VGND VGND VPWR VPWR net2041 sky130_fd_sc_hd__dlygate4sd3_1
X_11003_ net2282 net988 net341 VGND VGND VPWR VPWR _02747_ sky130_fd_sc_hd__mux2_1
XFILLER_120_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout870 _05540_ VGND VGND VPWR VPWR net870 sky130_fd_sc_hd__clkbuf_2
XFILLER_77_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout881 net882 VGND VGND VPWR VPWR net881 sky130_fd_sc_hd__buf_1
Xfanout892 _05528_ VGND VGND VPWR VPWR net892 sky130_fd_sc_hd__clkbuf_2
XFILLER_92_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12954_ clknet_leaf_207_clk _01648_ VGND VGND VPWR VPWR data_array.data0\[13\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_45_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1090 data_array.data1\[4\]\[21\] VGND VGND VPWR VPWR net2741 sky130_fd_sc_hd__dlygate4sd3_1
X_11905_ clknet_leaf_50_clk _00713_ VGND VGND VPWR VPWR data_array.data0\[5\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_193_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_193_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12885_ clknet_leaf_3_clk _01579_ VGND VGND VPWR VPWR data_array.data0\[12\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_178_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11836_ clknet_leaf_89_clk _00644_ VGND VGND VPWR VPWR data_array.data0\[7\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11767_ clknet_leaf_89_clk _00575_ VGND VGND VPWR VPWR data_array.data0\[8\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
X_13506_ clknet_leaf_36_clk _02135_ VGND VGND VPWR VPWR data_array.data1\[0\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_10718_ net1100 net2718 net490 VGND VGND VPWR VPWR _02463_ sky130_fd_sc_hd__mux2_1
X_14486_ clknet_leaf_161_clk _03109_ VGND VGND VPWR VPWR tag_array.dirty0\[5\] sky130_fd_sc_hd__dfxtp_1
X_11698_ clknet_leaf_231_clk _00506_ VGND VGND VPWR VPWR tag_array.tag1\[15\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13437_ clknet_leaf_238_clk _02067_ VGND VGND VPWR VPWR data_array.data1\[8\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload205 clknet_leaf_112_clk VGND VGND VPWR VPWR clkload205/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload216 clknet_leaf_123_clk VGND VGND VPWR VPWR clkload216/Y sky130_fd_sc_hd__clkinv_2
X_10649_ net2159 net865 net470 VGND VGND VPWR VPWR _02394_ sky130_fd_sc_hd__mux2_1
Xrebuffer2 fsm.tag_out0\[5\] VGND VGND VPWR VPWR net1653 sky130_fd_sc_hd__dlygate4sd1_1
Xclkload227 clknet_leaf_151_clk VGND VGND VPWR VPWR clkload227/Y sky130_fd_sc_hd__clkinv_2
Xclkload238 clknet_leaf_135_clk VGND VGND VPWR VPWR clkload238/Y sky130_fd_sc_hd__inv_6
XFILLER_173_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13368_ clknet_leaf_141_clk _01998_ VGND VGND VPWR VPWR tag_array.tag0\[2\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_77_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12319_ clknet_leaf_266_clk _00011_ VGND VGND VPWR VPWR data_array.rdata0\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13299_ clknet_leaf_16_clk _01929_ VGND VGND VPWR VPWR data_array.data0\[10\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2708 data_array.data1\[3\]\[35\] VGND VGND VPWR VPWR net4359 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2719 tag_array.tag0\[10\]\[6\] VGND VGND VPWR VPWR net4370 sky130_fd_sc_hd__dlygate4sd3_1
X_07860_ data_array.data1\[8\]\[38\] net1397 net1303 data_array.data1\[11\]\[38\]
+ _05062_ VGND VGND VPWR VPWR _05063_ sky130_fd_sc_hd__a221o_1
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06811_ net1614 _04103_ _04107_ net1188 VGND VGND VPWR VPWR _04110_ sky130_fd_sc_hd__a22o_1
XFILLER_110_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07791_ net1177 _04995_ _04999_ net1224 VGND VGND VPWR VPWR _05001_ sky130_fd_sc_hd__a22o_1
XFILLER_110_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06742_ data_array.data0\[8\]\[0\] net1367 net1273 data_array.data0\[11\]\[0\] _04046_
+ VGND VGND VPWR VPWR _04047_ sky130_fd_sc_hd__a221o_1
X_09530_ net709 net2305 net622 VGND VGND VPWR VPWR _01283_ sky130_fd_sc_hd__mux2_1
XFILLER_3_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09461_ net783 net3827 net651 VGND VGND VPWR VPWR _01214_ sky130_fd_sc_hd__mux2_1
X_06673_ tag_array.tag1\[5\]\[19\] net1576 net1480 tag_array.tag1\[6\]\[19\] VGND
+ VGND VPWR VPWR _03984_ sky130_fd_sc_hd__a22o_1
XFILLER_36_275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_184_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_184_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_24_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08412_ net139 net74 net1638 VGND VGND VPWR VPWR _05511_ sky130_fd_sc_hd__mux2_1
X_05624_ net164 VGND VGND VPWR VPWR _00189_ sky130_fd_sc_hd__inv_2
XFILLER_51_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09392_ net1099 net2608 net580 VGND VGND VPWR VPWR _01145_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_177_3770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08343_ net114 net49 net1643 VGND VGND VPWR VPWR _05465_ sky130_fd_sc_hd__mux2_1
XFILLER_149_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_3678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08274_ net99 net34 net1644 VGND VGND VPWR VPWR _05419_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_173_3689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07225_ data_array.data0\[13\]\[44\] net1586 net1490 data_array.data0\[14\]\[44\]
+ VGND VGND VPWR VPWR _04486_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_134_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07156_ data_array.data0\[8\]\[38\] net1396 net1302 data_array.data0\[11\]\[38\]
+ _04422_ VGND VGND VPWR VPWR _04423_ sky130_fd_sc_hd__a221o_1
XFILLER_152_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06107_ data_array.rdata0\[22\] net1135 net1112 data_array.rdata1\[22\] VGND VGND
+ VPWR VPWR net277 sky130_fd_sc_hd__a22o_1
XFILLER_145_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07087_ net1177 _04355_ _04359_ net1225 VGND VGND VPWR VPWR _04361_ sky130_fd_sc_hd__a22o_1
XFILLER_105_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06038_ fsm.tag_out0\[1\] net1120 _03482_ VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__a21o_1
XFILLER_105_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1109 _05420_ VGND VGND VPWR VPWR net1109 sky130_fd_sc_hd__buf_1
XFILLER_102_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07989_ net1226 _05175_ _05179_ net1178 VGND VGND VPWR VPWR _05181_ sky130_fd_sc_hd__a22o_1
X_09728_ net774 net2640 net678 VGND VGND VPWR VPWR _01480_ sky130_fd_sc_hd__mux2_1
XFILLER_41_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_175_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_175_clk
+ sky130_fd_sc_hd__clkbuf_8
X_09659_ net752 net3945 net613 VGND VGND VPWR VPWR _01411_ sky130_fd_sc_hd__mux2_1
XFILLER_42_223 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12670_ clknet_leaf_224_clk _01364_ VGND VGND VPWR VPWR data_array.data0\[15\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_151_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11621_ clknet_leaf_167_clk _00429_ VGND VGND VPWR VPWR tag_array.tag1\[3\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14340_ clknet_leaf_120_clk _02969_ VGND VGND VPWR VPWR data_array.data1\[11\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_13_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11552_ clknet_leaf_189_clk _00360_ VGND VGND VPWR VPWR tag_array.tag1\[6\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10503_ net932 net3537 net350 VGND VGND VPWR VPWR _02248_ sky130_fd_sc_hd__mux2_1
X_14271_ clknet_leaf_20_clk _02900_ VGND VGND VPWR VPWR data_array.data1\[12\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
X_11483_ clknet_leaf_152_clk _00292_ VGND VGND VPWR VPWR tag_array.valid0\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10434_ net2044 net918 net668 VGND VGND VPWR VPWR _02180_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13222_ clknet_leaf_52_clk _00118_ VGND VGND VPWR VPWR data_array.rdata1\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_143_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13153_ clknet_leaf_99_clk _01847_ VGND VGND VPWR VPWR tag_array.tag1\[8\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10365_ net738 net4152 net539 VGND VGND VPWR VPWR _02112_ sky130_fd_sc_hd__mux2_1
XFILLER_128_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12104_ clknet_leaf_245_clk _00912_ VGND VGND VPWR VPWR data_array.data1\[14\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
X_13084_ clknet_leaf_259_clk _01778_ VGND VGND VPWR VPWR data_array.data1\[13\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
X_10296_ net2413 net979 net640 VGND VGND VPWR VPWR _02043_ sky130_fd_sc_hd__mux2_1
XFILLER_78_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1610 net1612 VGND VGND VPWR VPWR net1610 sky130_fd_sc_hd__clkbuf_4
X_12035_ clknet_leaf_20_clk _00843_ VGND VGND VPWR VPWR data_array.data0\[6\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_72_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1621 net1624 VGND VGND VPWR VPWR net1621 sky130_fd_sc_hd__buf_4
Xfanout1632 _03506_ VGND VGND VPWR VPWR net1632 sky130_fd_sc_hd__buf_4
Xfanout1643 net1645 VGND VGND VPWR VPWR net1643 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13986_ clknet_leaf_256_clk _02615_ VGND VGND VPWR VPWR data_array.data1\[5\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_12937_ clknet_leaf_260_clk _01631_ VGND VGND VPWR VPWR data_array.data0\[13\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_166_clk clknet_5_24__leaf_clk VGND VGND VPWR VPWR clknet_leaf_166_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_61_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12868_ clknet_leaf_114_clk _01562_ VGND VGND VPWR VPWR data_array.data0\[12\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_138_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11819_ clknet_leaf_228_clk _00627_ VGND VGND VPWR VPWR data_array.data0\[7\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_12799_ clknet_leaf_141_clk _01493_ VGND VGND VPWR VPWR tag_array.tag1\[10\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_155_3342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14469_ clknet_leaf_5_clk _03092_ VGND VGND VPWR VPWR data_array.data1\[7\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
X_07010_ net1177 _04285_ _04289_ net1225 VGND VGND VPWR VPWR _04291_ sky130_fd_sc_hd__a22o_1
XFILLER_146_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08961_ net921 net2888 net431 VGND VGND VPWR VPWR _00717_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2505 tag_array.tag1\[7\]\[15\] VGND VGND VPWR VPWR net4156 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2516 tag_array.tag1\[14\]\[7\] VGND VGND VPWR VPWR net4167 sky130_fd_sc_hd__dlygate4sd3_1
X_07912_ net1179 _05105_ _05109_ net1227 VGND VGND VPWR VPWR _05111_ sky130_fd_sc_hd__a22o_1
Xhold2527 data_array.data0\[7\]\[30\] VGND VGND VPWR VPWR net4178 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2538 data_array.data0\[11\]\[8\] VGND VGND VPWR VPWR net4189 sky130_fd_sc_hd__dlygate4sd3_1
X_08892_ net936 net3909 net439 VGND VGND VPWR VPWR _00649_ sky130_fd_sc_hd__mux2_1
XFILLER_124_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1804 data_array.data1\[10\]\[49\] VGND VGND VPWR VPWR net3455 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2549 data_array.data0\[3\]\[57\] VGND VGND VPWR VPWR net4200 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1815 data_array.data1\[8\]\[38\] VGND VGND VPWR VPWR net3466 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07843_ data_array.data1\[1\]\[36\] net1604 net1508 data_array.data1\[2\]\[36\] VGND
+ VGND VPWR VPWR _05048_ sky130_fd_sc_hd__a22o_1
Xhold1826 tag_array.dirty1\[11\] VGND VGND VPWR VPWR net3477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1837 data_array.data1\[7\]\[15\] VGND VGND VPWR VPWR net3488 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_68_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1848 data_array.data1\[9\]\[61\] VGND VGND VPWR VPWR net3499 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1859 data_array.data0\[6\]\[55\] VGND VGND VPWR VPWR net3510 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07774_ data_array.data1\[4\]\[30\] net1393 net1299 data_array.data1\[7\]\[30\] _04984_
+ VGND VGND VPWR VPWR _04985_ sky130_fd_sc_hd__a221o_1
Xclone7 net852 VGND VGND VPWR VPWR net1658 sky130_fd_sc_hd__clkbuf_4
XFILLER_17_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09513_ net777 net4485 net621 VGND VGND VPWR VPWR _01266_ sky130_fd_sc_hd__mux2_1
XFILLER_140_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06725_ _04030_ _04031_ VGND VGND VPWR VPWR _00171_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_157_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_157_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_175_3718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06656_ tag_array.tag1\[0\]\[17\] net1418 net1324 tag_array.tag1\[3\]\[17\] _03968_
+ VGND VGND VPWR VPWR _03969_ sky130_fd_sc_hd__a221o_1
X_09444_ net891 net2599 net580 VGND VGND VPWR VPWR _01197_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_175_3729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_166_Right_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09375_ net902 net2679 net405 VGND VGND VPWR VPWR _01128_ sky130_fd_sc_hd__mux2_1
X_06587_ tag_array.tag1\[13\]\[11\] net1576 net1480 tag_array.tag1\[14\]\[11\] VGND
+ VGND VPWR VPWR _03906_ sky130_fd_sc_hd__a22o_1
X_08326_ net1125 _05453_ VGND VGND VPWR VPWR _05454_ sky130_fd_sc_hd__and2_1
XFILLER_71_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08257_ net1651 net1162 net21 VGND VGND VPWR VPWR _05406_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_31_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07208_ net1179 _04465_ _04469_ net1227 VGND VGND VPWR VPWR _04471_ sky130_fd_sc_hd__a22o_1
XFILLER_180_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08188_ _03320_ _03326_ _03327_ _03332_ fsm.state\[2\] VGND VGND VPWR VPWR _05358_
+ sky130_fd_sc_hd__o41a_1
XFILLER_106_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_104_Left_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07139_ data_array.data0\[1\]\[36\] net1601 net1505 data_array.data0\[2\]\[36\] VGND
+ VGND VPWR VPWR _04408_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_83_Right_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10150_ net945 net4033 net363 VGND VGND VPWR VPWR _01898_ sky130_fd_sc_hd__mux2_1
XFILLER_161_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput270 net270 VGND VGND VPWR VPWR mem_wdata[16] sky130_fd_sc_hd__buf_2
Xoutput281 net281 VGND VGND VPWR VPWR mem_wdata[26] sky130_fd_sc_hd__buf_2
Xoutput292 net292 VGND VGND VPWR VPWR mem_wdata[36] sky130_fd_sc_hd__buf_2
XFILLER_88_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10081_ net699 net4303 net600 VGND VGND VPWR VPWR _01830_ sky130_fd_sc_hd__mux2_1
XFILLER_0_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13840_ clknet_leaf_19_clk _02469_ VGND VGND VPWR VPWR data_array.data1\[3\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_113_Left_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13771_ clknet_leaf_36_clk _02400_ VGND VGND VPWR VPWR data_array.data1\[2\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_148_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_148_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10983_ net2440 net1068 net343 VGND VGND VPWR VPWR _02727_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_92_Right_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12722_ clknet_leaf_165_clk _01416_ VGND VGND VPWR VPWR tag_array.tag0\[7\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_133_Right_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12653_ clknet_leaf_241_clk _01347_ VGND VGND VPWR VPWR data_array.data0\[15\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
X_11604_ clknet_leaf_232_clk _00412_ VGND VGND VPWR VPWR tag_array.tag1\[4\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12584_ clknet_leaf_157_clk _01278_ VGND VGND VPWR VPWR tag_array.tag0\[10\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_96_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14323_ clknet_leaf_43_clk _02952_ VGND VGND VPWR VPWR data_array.data1\[11\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_129_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11535_ clknet_leaf_32_clk _00343_ VGND VGND VPWR VPWR tag_array.tag1\[6\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_183_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14254_ clknet_leaf_77_clk _02883_ VGND VGND VPWR VPWR data_array.data1\[12\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_150_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11466_ clknet_leaf_14_clk _00276_ VGND VGND VPWR VPWR data_array.data0\[0\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_139_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13205_ clknet_leaf_80_clk _00100_ VGND VGND VPWR VPWR data_array.rdata1\[42\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_74_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10417_ net1769 net984 net667 VGND VGND VPWR VPWR _02163_ sky130_fd_sc_hd__mux2_1
XFILLER_87_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11397_ clknet_leaf_33_clk _00207_ VGND VGND VPWR VPWR tag_array.tag1\[7\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_111_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14185_ clknet_leaf_91_clk _02814_ VGND VGND VPWR VPWR data_array.data0\[2\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_140_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13136_ clknet_leaf_127_clk _01830_ VGND VGND VPWR VPWR tag_array.tag0\[3\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_180_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10348_ net708 net2280 net593 VGND VGND VPWR VPWR _02095_ sky130_fd_sc_hd__mux2_1
XFILLER_124_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10279_ net2259 net1044 net637 VGND VGND VPWR VPWR _02026_ sky130_fd_sc_hd__mux2_1
X_13067_ clknet_leaf_46_clk _01761_ VGND VGND VPWR VPWR data_array.data1\[13\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout1440 net1447 VGND VGND VPWR VPWR net1440 sky130_fd_sc_hd__buf_2
XFILLER_38_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12018_ clknet_leaf_26_clk _00826_ VGND VGND VPWR VPWR data_array.data0\[6\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout1451 net1453 VGND VGND VPWR VPWR net1451 sky130_fd_sc_hd__clkbuf_4
Xfanout1462 net1464 VGND VGND VPWR VPWR net1462 sky130_fd_sc_hd__clkbuf_4
XFILLER_78_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1473 net1477 VGND VGND VPWR VPWR net1473 sky130_fd_sc_hd__clkbuf_2
Xfanout1484 net1486 VGND VGND VPWR VPWR net1484 sky130_fd_sc_hd__clkbuf_4
Xfanout1495 net1518 VGND VGND VPWR VPWR net1495 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_109_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1012 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13969_ clknet_leaf_57_clk _02598_ VGND VGND VPWR VPWR data_array.data1\[5\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_139_clk clknet_5_31__leaf_clk VGND VGND VPWR VPWR clknet_leaf_139_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_81_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06510_ tag_array.tag1\[13\]\[4\] net1552 net1456 tag_array.tag1\[14\]\[4\] VGND
+ VGND VPWR VPWR _03836_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07490_ data_array.data1\[12\]\[4\] net1393 net1299 data_array.data1\[15\]\[4\] _04726_
+ VGND VGND VPWR VPWR _04727_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_17_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06441_ tag_array.tag0\[8\]\[23\] net1409 net1315 tag_array.tag0\[11\]\[23\] _03772_
+ VGND VGND VPWR VPWR _03773_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_100_Right_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09160_ net901 net3831 net570 VGND VGND VPWR VPWR _00914_ sky130_fd_sc_hd__mux2_1
X_06372_ net1182 _03705_ _03709_ net1230 VGND VGND VPWR VPWR _03711_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_170_3626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08111_ _05290_ _05291_ VGND VGND VPWR VPWR _00120_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_170_3637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09091_ net921 net2354 net415 VGND VGND VPWR VPWR _00845_ sky130_fd_sc_hd__mux2_1
X_08042_ data_array.data1\[4\]\[54\] net1353 net1259 data_array.data1\[7\]\[54\] _05228_
+ VGND VGND VPWR VPWR _05229_ sky130_fd_sc_hd__a221o_1
XFILLER_31_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold901 data_array.data0\[11\]\[35\] VGND VGND VPWR VPWR net2552 sky130_fd_sc_hd__dlygate4sd3_1
Xhold912 tag_array.tag0\[13\]\[8\] VGND VGND VPWR VPWR net2563 sky130_fd_sc_hd__dlygate4sd3_1
Xhold923 data_array.data0\[2\]\[8\] VGND VGND VPWR VPWR net2574 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_843 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold934 data_array.data1\[12\]\[44\] VGND VGND VPWR VPWR net2585 sky130_fd_sc_hd__dlygate4sd3_1
Xhold945 data_array.data0\[13\]\[22\] VGND VGND VPWR VPWR net2596 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold956 tag_array.tag0\[0\]\[24\] VGND VGND VPWR VPWR net2607 sky130_fd_sc_hd__dlygate4sd3_1
Xhold967 data_array.data1\[12\]\[7\] VGND VGND VPWR VPWR net2618 sky130_fd_sc_hd__dlygate4sd3_1
Xhold978 tag_array.tag1\[15\]\[21\] VGND VGND VPWR VPWR net2629 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold989 tag_array.tag1\[10\]\[4\] VGND VGND VPWR VPWR net2640 sky130_fd_sc_hd__dlygate4sd3_1
X_09993_ net856 net3298 net372 VGND VGND VPWR VPWR _01742_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_168_3588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_3599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2302 tag_array.tag1\[10\]\[12\] VGND VGND VPWR VPWR net3953 sky130_fd_sc_hd__dlygate4sd3_1
X_08944_ net988 net2788 net430 VGND VGND VPWR VPWR _00700_ sky130_fd_sc_hd__mux2_1
Xhold2313 data_array.data0\[7\]\[56\] VGND VGND VPWR VPWR net3964 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2324 data_array.data0\[3\]\[24\] VGND VGND VPWR VPWR net3975 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2335 data_array.data1\[9\]\[22\] VGND VGND VPWR VPWR net3986 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2346 data_array.data0\[2\]\[1\] VGND VGND VPWR VPWR net3997 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1601 data_array.data1\[5\]\[42\] VGND VGND VPWR VPWR net3252 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1612 data_array.data0\[10\]\[13\] VGND VGND VPWR VPWR net3263 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2357 tag_array.tag0\[8\]\[20\] VGND VGND VPWR VPWR net4008 sky130_fd_sc_hd__dlygate4sd3_1
X_08875_ net1006 net2470 net436 VGND VGND VPWR VPWR _00632_ sky130_fd_sc_hd__mux2_1
Xhold1623 tag_array.tag0\[9\]\[1\] VGND VGND VPWR VPWR net3274 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2368 tag_array.tag1\[3\]\[4\] VGND VGND VPWR VPWR net4019 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_635 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1634 tag_array.tag1\[11\]\[18\] VGND VGND VPWR VPWR net3285 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2379 tag_array.tag0\[5\]\[21\] VGND VGND VPWR VPWR net4030 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1645 data_array.data1\[10\]\[1\] VGND VGND VPWR VPWR net3296 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1656 tag_array.tag1\[13\]\[16\] VGND VGND VPWR VPWR net3307 sky130_fd_sc_hd__dlygate4sd3_1
X_07826_ data_array.data1\[13\]\[35\] net1525 net1429 data_array.data1\[14\]\[35\]
+ VGND VGND VPWR VPWR _05032_ sky130_fd_sc_hd__a22o_1
Xhold1667 tag_array.tag0\[9\]\[20\] VGND VGND VPWR VPWR net3318 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1678 data_array.data0\[15\]\[42\] VGND VGND VPWR VPWR net3329 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1689 tag_array.tag0\[4\]\[16\] VGND VGND VPWR VPWR net3340 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07757_ net1620 _04963_ _04967_ net1194 VGND VGND VPWR VPWR _04970_ sky130_fd_sc_hd__a22o_1
XFILLER_84_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06708_ tag_array.tag1\[9\]\[22\] net1551 net1455 tag_array.tag1\[10\]\[22\] VGND
+ VGND VPWR VPWR _04016_ sky130_fd_sc_hd__a22o_1
X_07688_ data_array.data1\[12\]\[22\] net1346 net1252 data_array.data1\[15\]\[22\]
+ _04906_ VGND VGND VPWR VPWR _04907_ sky130_fd_sc_hd__a221o_1
XFILLER_80_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09427_ net958 net4078 net586 VGND VGND VPWR VPWR _01180_ sky130_fd_sc_hd__mux2_1
XFILLER_52_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06639_ tag_array.tag1\[12\]\[16\] net1417 net1323 tag_array.tag1\[15\]\[16\] _03952_
+ VGND VGND VPWR VPWR _03953_ sky130_fd_sc_hd__a221o_1
X_09358_ net970 net4371 net402 VGND VGND VPWR VPWR _01111_ sky130_fd_sc_hd__mux2_1
X_08309_ net2154 net1064 net692 VGND VGND VPWR VPWR _00232_ sky130_fd_sc_hd__mux2_1
XFILLER_139_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09289_ net725 net3047 net564 VGND VGND VPWR VPWR _01043_ sky130_fd_sc_hd__mux2_1
XFILLER_138_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11320_ net1014 net3049 net801 VGND VGND VPWR VPWR _03063_ sky130_fd_sc_hd__mux2_1
XFILLER_153_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11251_ net1024 net3379 net677 VGND VGND VPWR VPWR _02994_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10202_ net998 net3829 net355 VGND VGND VPWR VPWR _01949_ sky130_fd_sc_hd__mux2_1
XFILLER_122_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11182_ net1045 net4449 net652 VGND VGND VPWR VPWR _02925_ sky130_fd_sc_hd__mux2_1
XFILLER_134_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10133_ net1012 net4092 net366 VGND VGND VPWR VPWR _01881_ sky130_fd_sc_hd__mux2_1
XFILLER_133_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10064_ net768 net2806 net599 VGND VGND VPWR VPWR _01813_ sky130_fd_sc_hd__mux2_1
XFILLER_85_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_121_Left_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2880 data_array.data0\[7\]\[22\] VGND VGND VPWR VPWR net4531 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2891 data_array.data0\[13\]\[20\] VGND VGND VPWR VPWR net4542 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13823_ clknet_leaf_17_clk _02452_ VGND VGND VPWR VPWR data_array.data1\[2\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13754_ clknet_leaf_246_clk _02383_ VGND VGND VPWR VPWR data_array.data1\[1\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_67_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10966_ net878 net3791 net529 VGND VGND VPWR VPWR _02711_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12705_ clknet_leaf_143_clk _01399_ VGND VGND VPWR VPWR tag_array.tag0\[8\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_71_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13685_ clknet_leaf_28_clk _02314_ VGND VGND VPWR VPWR data_array.data1\[15\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
X_10897_ net898 net2728 net518 VGND VGND VPWR VPWR _02642_ sky130_fd_sc_hd__mux2_1
XFILLER_148_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12636_ clknet_leaf_15_clk _01330_ VGND VGND VPWR VPWR data_array.data0\[15\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_100_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_130_Left_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12567_ clknet_leaf_185_clk _01261_ VGND VGND VPWR VPWR tag_array.tag0\[11\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_129_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14306_ clknet_leaf_259_clk _02935_ VGND VGND VPWR VPWR data_array.data1\[11\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11518_ clknet_leaf_129_clk _00326_ VGND VGND VPWR VPWR tag_array.tag1\[9\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12498_ clknet_leaf_242_clk _01192_ VGND VGND VPWR VPWR data_array.data1\[9\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold208 data_array.data1\[0\]\[34\] VGND VGND VPWR VPWR net1859 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold219 data_array.data1\[8\]\[32\] VGND VGND VPWR VPWR net1870 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14237_ clknet_leaf_229_clk _02866_ VGND VGND VPWR VPWR data_array.data1\[12\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_11449_ clknet_leaf_88_clk _00259_ VGND VGND VPWR VPWR data_array.data0\[0\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
X_14168_ clknet_leaf_222_clk _02797_ VGND VGND VPWR VPWR data_array.data0\[2\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_98_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13119_ clknet_leaf_180_clk _01813_ VGND VGND VPWR VPWR tag_array.tag0\[3\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_140_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06990_ data_array.data0\[13\]\[23\] net1561 net1465 data_array.data0\[14\]\[23\]
+ VGND VGND VPWR VPWR _04272_ sky130_fd_sc_hd__a22o_1
X_14099_ clknet_leaf_43_clk _02728_ VGND VGND VPWR VPWR data_array.data0\[1\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_85_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05941_ net128 net1157 _03420_ _03421_ VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__a22o_1
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1270 net1282 VGND VGND VPWR VPWR net1270 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_163_3496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05872_ net103 net1152 _03374_ _03375_ VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__a22o_1
Xfanout1281 net1282 VGND VGND VPWR VPWR net1281 sky130_fd_sc_hd__buf_2
X_08660_ net782 net4342 net495 VGND VGND VPWR VPWR _00419_ sky130_fd_sc_hd__mux2_1
XFILLER_27_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1292 net1293 VGND VGND VPWR VPWR net1292 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_1_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07611_ data_array.data1\[12\]\[15\] net1391 net1297 data_array.data1\[15\]\[15\]
+ _04836_ VGND VGND VPWR VPWR _04837_ sky130_fd_sc_hd__a221o_1
XFILLER_54_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08591_ net759 net4237 net536 VGND VGND VPWR VPWR _00350_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_124_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07542_ data_array.data1\[5\]\[9\] net1580 net1484 data_array.data1\[6\]\[9\] VGND
+ VGND VPWR VPWR _04774_ sky130_fd_sc_hd__a22o_1
Xclkbuf_5_22__f_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_5_22__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_81_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07473_ _04710_ _04711_ VGND VGND VPWR VPWR _00086_ sky130_fd_sc_hd__or2_1
X_09212_ net733 net3772 net630 VGND VGND VPWR VPWR _00966_ sky130_fd_sc_hd__mux2_1
X_06424_ tag_array.tag0\[1\]\[21\] net1598 net1502 tag_array.tag0\[2\]\[21\] VGND
+ VGND VPWR VPWR _03758_ sky130_fd_sc_hd__a22o_1
XFILLER_179_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09143_ net969 net3509 net566 VGND VGND VPWR VPWR _00897_ sky130_fd_sc_hd__mux2_1
X_06355_ tag_array.tag0\[0\]\[15\] net1402 net1308 tag_array.tag0\[3\]\[15\] _03694_
+ VGND VGND VPWR VPWR _03695_ sky130_fd_sc_hd__a221o_1
XFILLER_148_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09074_ net988 net4205 net414 VGND VGND VPWR VPWR _00828_ sky130_fd_sc_hd__mux2_1
XFILLER_147_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06286_ tag_array.tag0\[13\]\[9\] net1599 net1503 tag_array.tag0\[14\]\[9\] VGND
+ VGND VPWR VPWR _03632_ sky130_fd_sc_hd__a22o_1
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08025_ data_array.data1\[8\]\[53\] net1334 net1240 data_array.data1\[11\]\[53\]
+ _05212_ VGND VGND VPWR VPWR _05213_ sky130_fd_sc_hd__a221o_1
XFILLER_116_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold720 data_array.data0\[2\]\[54\] VGND VGND VPWR VPWR net2371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold731 data_array.data0\[4\]\[61\] VGND VGND VPWR VPWR net2382 sky130_fd_sc_hd__dlygate4sd3_1
Xhold742 tag_array.tag0\[11\]\[13\] VGND VGND VPWR VPWR net2393 sky130_fd_sc_hd__dlygate4sd3_1
Xhold753 data_array.data0\[1\]\[54\] VGND VGND VPWR VPWR net2404 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold764 tag_array.tag1\[14\]\[13\] VGND VGND VPWR VPWR net2415 sky130_fd_sc_hd__dlygate4sd3_1
Xhold775 data_array.data1\[3\]\[36\] VGND VGND VPWR VPWR net2426 sky130_fd_sc_hd__dlygate4sd3_1
Xhold786 tag_array.tag0\[4\]\[14\] VGND VGND VPWR VPWR net2437 sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 data_array.data1\[2\]\[60\] VGND VGND VPWR VPWR net2448 sky130_fd_sc_hd__dlygate4sd3_1
X_09976_ net926 net3822 net370 VGND VGND VPWR VPWR _01725_ sky130_fd_sc_hd__mux2_1
Xhold2110 tag_array.tag0\[6\]\[10\] VGND VGND VPWR VPWR net3761 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2121 tag_array.tag0\[13\]\[15\] VGND VGND VPWR VPWR net3772 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2132 data_array.data0\[14\]\[4\] VGND VGND VPWR VPWR net3783 sky130_fd_sc_hd__dlygate4sd3_1
X_08927_ net1058 net3797 net428 VGND VGND VPWR VPWR _00683_ sky130_fd_sc_hd__mux2_1
Xhold2143 data_array.data0\[9\]\[4\] VGND VGND VPWR VPWR net3794 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2154 tag_array.tag0\[8\]\[9\] VGND VGND VPWR VPWR net3805 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2165 data_array.data1\[10\]\[17\] VGND VGND VPWR VPWR net3816 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1420 tag_array.tag0\[9\]\[9\] VGND VGND VPWR VPWR net3071 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1431 data_array.data0\[0\]\[34\] VGND VGND VPWR VPWR net3082 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2176 tag_array.tag1\[11\]\[2\] VGND VGND VPWR VPWR net3827 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1442 data_array.data0\[9\]\[42\] VGND VGND VPWR VPWR net3093 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2187 data_array.data0\[6\]\[50\] VGND VGND VPWR VPWR net3838 sky130_fd_sc_hd__dlygate4sd3_1
X_08858_ net1072 net3730 net438 VGND VGND VPWR VPWR _00615_ sky130_fd_sc_hd__mux2_1
Xhold2198 data_array.data1\[7\]\[30\] VGND VGND VPWR VPWR net3849 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1453 tag_array.tag0\[2\]\[4\] VGND VGND VPWR VPWR net3104 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1464 data_array.data1\[13\]\[29\] VGND VGND VPWR VPWR net3115 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1475 data_array.data0\[12\]\[49\] VGND VGND VPWR VPWR net3126 sky130_fd_sc_hd__dlygate4sd3_1
X_07809_ data_array.data1\[8\]\[33\] net1398 net1304 data_array.data1\[11\]\[33\]
+ _05016_ VGND VGND VPWR VPWR _05017_ sky130_fd_sc_hd__a221o_1
Xhold1486 data_array.data1\[9\]\[58\] VGND VGND VPWR VPWR net3137 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1497 data_array.data1\[3\]\[57\] VGND VGND VPWR VPWR net3148 sky130_fd_sc_hd__dlygate4sd3_1
X_08789_ net1754 net1089 net444 VGND VGND VPWR VPWR _00547_ sky130_fd_sc_hd__mux2_1
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10820_ net1975 net950 net510 VGND VGND VPWR VPWR _02565_ sky130_fd_sc_hd__mux2_1
XFILLER_26_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10751_ net968 net4359 net491 VGND VGND VPWR VPWR _02496_ sky130_fd_sc_hd__mux2_1
XFILLER_38_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1079 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13470_ clknet_leaf_163_clk _02100_ VGND VGND VPWR VPWR tag_array.tag0\[15\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_10682_ net1914 net990 net484 VGND VGND VPWR VPWR _02427_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12421_ clknet_leaf_235_clk _01115_ VGND VGND VPWR VPWR data_array.data0\[14\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_127_916 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12352_ clknet_leaf_11_clk _00027_ VGND VGND VPWR VPWR data_array.rdata0\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11303_ net1082 net4323 net801 VGND VGND VPWR VPWR _03046_ sky130_fd_sc_hd__mux2_1
X_12283_ clknet_leaf_100_clk _01041_ VGND VGND VPWR VPWR tag_array.tag1\[13\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_153_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14022_ clknet_leaf_124_clk _02651_ VGND VGND VPWR VPWR data_array.data1\[5\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11234_ net1095 net4161 net681 VGND VGND VPWR VPWR _02977_ sky130_fd_sc_hd__mux2_1
XFILLER_4_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1025 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11165_ net858 net3729 net545 VGND VGND VPWR VPWR _02908_ sky130_fd_sc_hd__mux2_1
XFILLER_150_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10116_ net1081 net4315 net368 VGND VGND VPWR VPWR _01864_ sky130_fd_sc_hd__mux2_1
X_11096_ net2014 net876 net330 VGND VGND VPWR VPWR _02839_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_145_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10047_ net899 net3636 net554 VGND VGND VPWR VPWR _01796_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_69_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold80 data_array.data1\[2\]\[19\] VGND VGND VPWR VPWR net1731 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold91 data_array.data1\[0\]\[19\] VGND VGND VPWR VPWR net1742 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_64_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_106_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13806_ clknet_leaf_74_clk _02435_ VGND VGND VPWR VPWR data_array.data1\[2\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11998_ clknet_leaf_14_clk _00806_ VGND VGND VPWR VPWR data_array.data0\[6\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13737_ clknet_leaf_73_clk _02366_ VGND VGND VPWR VPWR data_array.data1\[1\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_82_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10949_ net944 net3767 net526 VGND VGND VPWR VPWR _02694_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_82_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_70_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_70_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_177_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13668_ clknet_leaf_30_clk _02297_ VGND VGND VPWR VPWR data_array.data1\[15\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_176_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12619_ clknet_leaf_261_clk _01313_ VGND VGND VPWR VPWR data_array.data0\[15\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13599_ clknet_leaf_92_clk _02228_ VGND VGND VPWR VPWR data_array.data0\[9\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_129_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06140_ data_array.rdata0\[55\] net1138 net1113 data_array.rdata1\[55\] VGND VGND
+ VPWR VPWR net313 sky130_fd_sc_hd__a22o_1
XFILLER_157_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06071_ net1159 net18 fsm.tag_out1\[18\] net1133 VGND VGND VPWR VPWR _03499_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_165_3525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_3536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09830_ net889 net3382 net387 VGND VGND VPWR VPWR _01581_ sky130_fd_sc_hd__mux2_1
Xfanout507 net512 VGND VGND VPWR VPWR net507 sky130_fd_sc_hd__buf_4
Xfanout518 _05599_ VGND VGND VPWR VPWR net518 sky130_fd_sc_hd__clkbuf_8
Xfanout529 net530 VGND VGND VPWR VPWR net529 sky130_fd_sc_hd__clkbuf_8
XFILLER_112_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_182_3850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_3861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09761_ net2370 net742 net672 VGND VGND VPWR VPWR _01513_ sky130_fd_sc_hd__mux2_1
X_06973_ data_array.data0\[12\]\[21\] net1366 net1272 data_array.data0\[15\]\[21\]
+ _04256_ VGND VGND VPWR VPWR _04257_ sky130_fd_sc_hd__a221o_1
XFILLER_100_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08712_ net2547 net775 net469 VGND VGND VPWR VPWR _00471_ sky130_fd_sc_hd__mux2_1
X_05924_ net851 data_array.rdata0\[31\] net1148 VGND VGND VPWR VPWR _03410_ sky130_fd_sc_hd__o21a_1
X_09692_ net720 net3315 net605 VGND VGND VPWR VPWR _01444_ sky130_fd_sc_hd__mux2_1
XFILLER_55_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08643_ net1795 net750 net511 VGND VGND VPWR VPWR _00402_ sky130_fd_sc_hd__mux2_1
X_05855_ data_array.rdata0\[8\] net847 net1143 VGND VGND VPWR VPWR _03364_ sky130_fd_sc_hd__o21a_1
XFILLER_82_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08574_ _05352_ net812 VGND VGND VPWR VPWR _05602_ sky130_fd_sc_hd__and2_1
XFILLER_81_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_05786_ _03295_ _03297_ _03299_ _03302_ VGND VGND VPWR VPWR _03303_ sky130_fd_sc_hd__or4_1
X_07525_ data_array.data1\[4\]\[7\] net1399 net1305 data_array.data1\[7\]\[7\] _04758_
+ VGND VGND VPWR VPWR _04759_ sky130_fd_sc_hd__a221o_1
XFILLER_168_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_61_clk clknet_5_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_61_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_34_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07456_ data_array.data1\[9\]\[1\] net1520 net1424 data_array.data1\[10\]\[1\] VGND
+ VGND VPWR VPWR _04696_ sky130_fd_sc_hd__a22o_1
X_06407_ tag_array.tag0\[13\]\[20\] net1560 net1464 tag_array.tag0\[14\]\[20\] VGND
+ VGND VPWR VPWR _03742_ sky130_fd_sc_hd__a22o_1
XFILLER_41_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07387_ data_array.data0\[8\]\[59\] net1379 net1285 data_array.data0\[11\]\[59\]
+ _04632_ VGND VGND VPWR VPWR _04633_ sky130_fd_sc_hd__a221o_1
XFILLER_182_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09126_ net1038 net3731 net568 VGND VGND VPWR VPWR _00880_ sky130_fd_sc_hd__mux2_1
XFILLER_176_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06338_ net1637 _03673_ _03677_ net1211 VGND VGND VPWR VPWR _03680_ sky130_fd_sc_hd__a22o_1
XFILLER_175_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09057_ net1058 net3092 net412 VGND VGND VPWR VPWR _00811_ sky130_fd_sc_hd__mux2_1
X_06269_ tag_array.tag0\[12\]\[7\] net1409 net1315 tag_array.tag0\[15\]\[7\] _03616_
+ VGND VGND VPWR VPWR _03617_ sky130_fd_sc_hd__a221o_1
XFILLER_135_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08008_ data_array.data1\[1\]\[51\] net1522 net1426 data_array.data1\[2\]\[51\] VGND
+ VGND VPWR VPWR _05198_ sky130_fd_sc_hd__a22o_1
Xhold550 data_array.data1\[2\]\[23\] VGND VGND VPWR VPWR net2201 sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 data_array.data1\[4\]\[8\] VGND VGND VPWR VPWR net2212 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold572 data_array.data1\[2\]\[13\] VGND VGND VPWR VPWR net2223 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold583 data_array.data0\[1\]\[37\] VGND VGND VPWR VPWR net2234 sky130_fd_sc_hd__dlygate4sd3_1
Xhold594 data_array.data1\[8\]\[39\] VGND VGND VPWR VPWR net2245 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_173_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_538 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09959_ net992 net2477 net375 VGND VGND VPWR VPWR _01708_ sky130_fd_sc_hd__mux2_1
XFILLER_66_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_86_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12970_ clknet_leaf_107_clk _01664_ VGND VGND VPWR VPWR tag_array.tag0\[4\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_181_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1250 tag_array.dirty0\[10\] VGND VGND VPWR VPWR net2901 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1261 data_array.data1\[2\]\[42\] VGND VGND VPWR VPWR net2912 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11921_ clknet_leaf_52_clk _00729_ VGND VGND VPWR VPWR data_array.data0\[5\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1272 data_array.data0\[3\]\[61\] VGND VGND VPWR VPWR net2923 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1283 data_array.data0\[10\]\[20\] VGND VGND VPWR VPWR net2934 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1294 data_array.data0\[11\]\[20\] VGND VGND VPWR VPWR net2945 sky130_fd_sc_hd__dlygate4sd3_1
X_11852_ clknet_leaf_221_clk _00660_ VGND VGND VPWR VPWR data_array.data0\[7\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_122_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10803_ net1838 net1016 net505 VGND VGND VPWR VPWR _02548_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ clknet_leaf_61_clk _00591_ VGND VGND VPWR VPWR data_array.data0\[8\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_52_clk clknet_5_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_52_clk sky130_fd_sc_hd__clkbuf_8
X_13522_ clknet_leaf_66_clk _02151_ VGND VGND VPWR VPWR data_array.data1\[0\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_24_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10734_ net1038 net4234 net496 VGND VGND VPWR VPWR _02479_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_24_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13453_ clknet_leaf_160_clk _02083_ VGND VGND VPWR VPWR tag_array.tag0\[1\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_10665_ net2223 net1056 net481 VGND VGND VPWR VPWR _02410_ sky130_fd_sc_hd__mux2_1
XFILLER_167_882 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12404_ clknet_leaf_22_clk _01098_ VGND VGND VPWR VPWR data_array.data0\[14\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_13384_ clknet_leaf_68_clk _02014_ VGND VGND VPWR VPWR data_array.data1\[8\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_10596_ net1957 net1078 net467 VGND VGND VPWR VPWR _02341_ sky130_fd_sc_hd__mux2_1
XFILLER_12_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12335_ clknet_leaf_253_clk _00008_ VGND VGND VPWR VPWR data_array.rdata0\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_182_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12266_ clknet_leaf_130_clk _01024_ VGND VGND VPWR VPWR tag_array.tag1\[14\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_108_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_147_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14005_ clknet_leaf_25_clk _02634_ VGND VGND VPWR VPWR data_array.data1\[5\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
X_11217_ net907 net4536 net648 VGND VGND VPWR VPWR _02960_ sky130_fd_sc_hd__mux2_1
X_12197_ clknet_leaf_182_clk _00150_ VGND VGND VPWR VPWR fsm.tag_out0\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_1_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11148_ net924 net4242 net541 VGND VGND VPWR VPWR _02891_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_143_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_143_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_160_3433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11079_ net3232 net946 net328 VGND VGND VPWR VPWR _02822_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_160_3444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05640_ net18 fsm.tag_out0\[18\] VGND VGND VPWR VPWR _03157_ sky130_fd_sc_hd__xor2_1
XFILLER_17_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_43_clk clknet_5_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_43_clk sky130_fd_sc_hd__clkbuf_8
X_07310_ data_array.data0\[12\]\[52\] net1357 net1263 data_array.data0\[15\]\[52\]
+ _04562_ VGND VGND VPWR VPWR _04563_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_22_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08290_ net1126 _05429_ VGND VGND VPWR VPWR _05430_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_158_3395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07241_ net1216 _04495_ _04499_ net1168 VGND VGND VPWR VPWR _04501_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_119_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07172_ data_array.data0\[5\]\[39\] net1538 net1442 data_array.data0\[6\]\[39\] VGND
+ VGND VPWR VPWR _04438_ sky130_fd_sc_hd__a22o_1
X_06123_ data_array.rdata0\[38\] net1139 net1115 data_array.rdata1\[38\] VGND VGND
+ VPWR VPWR net294 sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_136_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06054_ fsm.tag_out0\[9\] net1121 _03490_ VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_184_3901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_184_3912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_180_3809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09813_ net957 net4184 net390 VGND VGND VPWR VPWR _01564_ sky130_fd_sc_hd__mux2_1
Xfanout337 net340 VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__buf_4
XFILLER_59_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout348 net350 VGND VGND VPWR VPWR net348 sky130_fd_sc_hd__buf_4
XFILLER_98_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout359 net360 VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__buf_4
X_09744_ net710 net4151 net675 VGND VGND VPWR VPWR _01496_ sky130_fd_sc_hd__mux2_1
XFILLER_101_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06956_ _04240_ _04241_ VGND VGND VPWR VPWR _00010_ sky130_fd_sc_hd__or2_1
XFILLER_28_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_05907_ data_array.rdata1\[25\] net828 net837 VGND VGND VPWR VPWR _03399_ sky130_fd_sc_hd__a21o_1
X_09675_ net789 net3670 net605 VGND VGND VPWR VPWR _01427_ sky130_fd_sc_hd__mux2_1
X_06887_ data_array.data0\[4\]\[13\] net1361 net1267 data_array.data0\[7\]\[13\] _04178_
+ VGND VGND VPWR VPWR _04179_ sky130_fd_sc_hd__a221o_1
X_08626_ net719 net2517 net517 VGND VGND VPWR VPWR _00385_ sky130_fd_sc_hd__mux2_1
X_05838_ data_array.rdata1\[2\] net830 net839 VGND VGND VPWR VPWR _03353_ sky130_fd_sc_hd__a21o_1
X_08557_ net728 net3201 net588 VGND VGND VPWR VPWR _00325_ sky130_fd_sc_hd__mux2_1
XFILLER_74_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05769_ net20 fsm.tag_out1\[20\] VGND VGND VPWR VPWR _03286_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_34_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_34_clk sky130_fd_sc_hd__clkbuf_8
X_07508_ data_array.data1\[8\]\[6\] net1329 net1235 data_array.data1\[11\]\[6\] _04742_
+ VGND VGND VPWR VPWR _04743_ sky130_fd_sc_hd__a221o_1
XFILLER_74_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08488_ _03514_ _03523_ net825 VGND VGND VPWR VPWR _05562_ sky130_fd_sc_hd__or3_1
XFILLER_11_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07439_ net1170 _04675_ _04679_ net1218 VGND VGND VPWR VPWR _04681_ sky130_fd_sc_hd__a22o_1
XFILLER_50_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10450_ net352 net4458 net800 VGND VGND VPWR VPWR _02196_ sky130_fd_sc_hd__mux2_1
XFILLER_6_328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09109_ net1106 net4491 net566 VGND VGND VPWR VPWR _00863_ sky130_fd_sc_hd__mux2_1
XFILLER_108_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10381_ net353 net3918 net544 VGND VGND VPWR VPWR _02127_ sky130_fd_sc_hd__mux2_1
X_12120_ clknet_leaf_171_clk _00928_ VGND VGND VPWR VPWR tag_array.tag0\[12\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12051_ clknet_leaf_207_clk _00859_ VGND VGND VPWR VPWR data_array.data0\[6\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold380 data_array.data1\[8\]\[5\] VGND VGND VPWR VPWR net2031 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold391 tag_array.tag1\[2\]\[3\] VGND VGND VPWR VPWR net2042 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11002_ net2481 net992 net341 VGND VGND VPWR VPWR _02746_ sky130_fd_sc_hd__mux2_1
XFILLER_77_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout860 _05544_ VGND VGND VPWR VPWR net860 sky130_fd_sc_hd__clkbuf_2
Xfanout871 _05540_ VGND VGND VPWR VPWR net871 sky130_fd_sc_hd__clkbuf_1
Xfanout882 _05534_ VGND VGND VPWR VPWR net882 sky130_fd_sc_hd__clkbuf_2
XFILLER_120_988 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout893 _05528_ VGND VGND VPWR VPWR net893 sky130_fd_sc_hd__clkbuf_1
XFILLER_92_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12953_ clknet_leaf_234_clk _01647_ VGND VGND VPWR VPWR data_array.data0\[13\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_133_83 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1080 tag_array.tag0\[10\]\[24\] VGND VGND VPWR VPWR net2731 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1091 data_array.data0\[0\]\[37\] VGND VGND VPWR VPWR net2742 sky130_fd_sc_hd__dlygate4sd3_1
X_11904_ clknet_leaf_93_clk _00712_ VGND VGND VPWR VPWR data_array.data0\[5\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_46_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12884_ clknet_leaf_224_clk _01578_ VGND VGND VPWR VPWR data_array.data0\[12\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
X_11835_ clknet_leaf_217_clk _00643_ VGND VGND VPWR VPWR data_array.data0\[7\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_25_clk clknet_5_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_8
X_11766_ clknet_leaf_260_clk _00574_ VGND VGND VPWR VPWR data_array.data0\[8\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_158_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13505_ clknet_leaf_252_clk _02134_ VGND VGND VPWR VPWR data_array.data1\[0\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_10717_ net1104 net4489 net490 VGND VGND VPWR VPWR _02462_ sky130_fd_sc_hd__mux2_1
X_14485_ clknet_leaf_161_clk _03108_ VGND VGND VPWR VPWR tag_array.dirty0\[4\] sky130_fd_sc_hd__dfxtp_1
X_11697_ clknet_leaf_134_clk _00505_ VGND VGND VPWR VPWR tag_array.tag1\[15\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13436_ clknet_leaf_22_clk _02066_ VGND VGND VPWR VPWR data_array.data1\[8\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
X_10648_ net1736 net870 net475 VGND VGND VPWR VPWR _02393_ sky130_fd_sc_hd__mux2_1
XFILLER_9_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload206 clknet_leaf_113_clk VGND VGND VPWR VPWR clkload206/Y sky130_fd_sc_hd__inv_6
XFILLER_167_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload217 clknet_leaf_124_clk VGND VGND VPWR VPWR clkload217/Y sky130_fd_sc_hd__clkinv_4
Xrebuffer3 _03207_ VGND VGND VPWR VPWR net1654 sky130_fd_sc_hd__dlygate4sd1_1
Xclkload228 clknet_leaf_152_clk VGND VGND VPWR VPWR clkload228/Y sky130_fd_sc_hd__inv_8
Xclkload239 clknet_leaf_136_clk VGND VGND VPWR VPWR clkload239/Y sky130_fd_sc_hd__clkinvlp_4
X_13367_ clknet_leaf_163_clk _01997_ VGND VGND VPWR VPWR tag_array.tag0\[2\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_154_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10579_ net891 net3096 net455 VGND VGND VPWR VPWR _02324_ sky130_fd_sc_hd__mux2_1
XFILLER_154_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12318_ clknet_leaf_185_clk _00000_ VGND VGND VPWR VPWR data_array.rdata0\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_77_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_844 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13298_ clknet_leaf_94_clk _01928_ VGND VGND VPWR VPWR data_array.data0\[10\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_170_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12249_ clknet_leaf_195_clk _01007_ VGND VGND VPWR VPWR tag_array.tag1\[14\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2709 tag_array.tag1\[5\]\[20\] VGND VGND VPWR VPWR net4360 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06810_ data_array.data0\[4\]\[6\] net1331 net1237 data_array.data0\[7\]\[6\] _04108_
+ VGND VGND VPWR VPWR _04109_ sky130_fd_sc_hd__a221o_1
XFILLER_95_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07790_ net1203 _04993_ _04997_ net1628 VGND VGND VPWR VPWR _05000_ sky130_fd_sc_hd__a22o_1
XFILLER_3_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_147_Right_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06741_ data_array.data0\[9\]\[0\] net1555 net1459 data_array.data0\[10\]\[0\] VGND
+ VGND VPWR VPWR _04046_ sky130_fd_sc_hd__a22o_1
XFILLER_97_1043 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09460_ net786 net4160 net650 VGND VGND VPWR VPWR _01213_ sky130_fd_sc_hd__mux2_1
XFILLER_97_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06672_ tag_array.tag1\[8\]\[19\] net1404 net1310 tag_array.tag1\[11\]\[19\] _03982_
+ VGND VGND VPWR VPWR _03983_ sky130_fd_sc_hd__a221o_1
XFILLER_36_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08411_ net2297 net928 net687 VGND VGND VPWR VPWR _00266_ sky130_fd_sc_hd__mux2_1
X_05623_ fsm.tag_out0\[18\] VGND VGND VPWR VPWR _03145_ sky130_fd_sc_hd__inv_2
X_09391_ net1101 net2988 net579 VGND VGND VPWR VPWR _01144_ sky130_fd_sc_hd__mux2_1
XFILLER_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_177_3760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_16_clk clknet_5_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_8
X_08342_ net1929 net1020 net687 VGND VGND VPWR VPWR _00243_ sky130_fd_sc_hd__mux2_1
XFILLER_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08273_ net1161 fsm.state\[2\] VGND VGND VPWR VPWR _05418_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_173_3679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07224_ data_array.data0\[0\]\[44\] net1395 net1301 data_array.data0\[3\]\[44\] _04484_
+ VGND VGND VPWR VPWR _04485_ sky130_fd_sc_hd__a221o_1
XFILLER_34_1071 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07155_ data_array.data0\[9\]\[38\] net1585 net1489 data_array.data0\[10\]\[38\]
+ VGND VGND VPWR VPWR _04422_ sky130_fd_sc_hd__a22o_1
XFILLER_106_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06106_ data_array.rdata0\[21\] net1136 net1117 data_array.rdata1\[21\] VGND VGND
+ VPWR VPWR net276 sky130_fd_sc_hd__a22o_1
XFILLER_133_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07086_ net1203 _04353_ _04357_ net1629 VGND VGND VPWR VPWR _04360_ sky130_fd_sc_hd__a22o_1
XFILLER_65_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06037_ net1158 net31 fsm.tag_out1\[1\] net1133 VGND VGND VPWR VPWR _03482_ sky130_fd_sc_hd__a22o_1
XFILLER_160_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07988_ net1203 _05173_ _05177_ net1629 VGND VGND VPWR VPWR _05180_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_114_Right_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09727_ net779 net4585 net677 VGND VGND VPWR VPWR _01479_ sky130_fd_sc_hd__mux2_1
XFILLER_28_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06939_ data_array.data0\[13\]\[18\] net1534 net1438 data_array.data0\[14\]\[18\]
+ VGND VGND VPWR VPWR _04226_ sky130_fd_sc_hd__a22o_1
XFILLER_27_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09658_ net754 net3010 net613 VGND VGND VPWR VPWR _01410_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08609_ net786 net4355 net525 VGND VGND VPWR VPWR _00368_ sky130_fd_sc_hd__mux2_1
XFILLER_82_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09589_ net993 net3848 net399 VGND VGND VPWR VPWR _01341_ sky130_fd_sc_hd__mux2_1
X_11620_ clknet_leaf_33_clk _00428_ VGND VGND VPWR VPWR tag_array.tag1\[3\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_179_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11551_ clknet_leaf_127_clk _00359_ VGND VGND VPWR VPWR tag_array.tag1\[6\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10502_ net939 net3615 net348 VGND VGND VPWR VPWR _02247_ sky130_fd_sc_hd__mux2_1
X_14270_ clknet_leaf_216_clk _02899_ VGND VGND VPWR VPWR data_array.data1\[12\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_98_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11482_ clknet_leaf_174_clk _00291_ VGND VGND VPWR VPWR tag_array.valid1\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_109_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13221_ clknet_leaf_211_clk _00117_ VGND VGND VPWR VPWR data_array.rdata1\[58\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_59_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10433_ net2229 net922 net669 VGND VGND VPWR VPWR _02179_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13152_ clknet_leaf_168_clk _01846_ VGND VGND VPWR VPWR tag_array.tag1\[8\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_88_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10364_ net744 net2689 net538 VGND VGND VPWR VPWR _02111_ sky130_fd_sc_hd__mux2_1
X_12103_ clknet_leaf_56_clk _00911_ VGND VGND VPWR VPWR data_array.data1\[14\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
X_13083_ clknet_leaf_8_clk _01777_ VGND VGND VPWR VPWR data_array.data1\[13\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
X_10295_ net1870 net981 net633 VGND VGND VPWR VPWR _02042_ sky130_fd_sc_hd__mux2_1
XFILLER_105_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1600 net1613 VGND VGND VPWR VPWR net1600 sky130_fd_sc_hd__clkbuf_2
X_12034_ clknet_leaf_87_clk _00842_ VGND VGND VPWR VPWR data_array.data0\[6\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout1611 net1612 VGND VGND VPWR VPWR net1611 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_72_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1622 net1624 VGND VGND VPWR VPWR net1622 sky130_fd_sc_hd__buf_4
Xfanout1633 net1634 VGND VGND VPWR VPWR net1633 sky130_fd_sc_hd__buf_4
Xfanout1644 net1645 VGND VGND VPWR VPWR net1644 sky130_fd_sc_hd__buf_4
XFILLER_78_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout690 _05417_ VGND VGND VPWR VPWR net690 sky130_fd_sc_hd__clkbuf_4
X_13985_ clknet_leaf_269_clk _02614_ VGND VGND VPWR VPWR data_array.data1\[5\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_5_3__f_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_5_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_12936_ clknet_leaf_124_clk _01630_ VGND VGND VPWR VPWR data_array.data0\[13\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12867_ clknet_leaf_242_clk _01561_ VGND VGND VPWR VPWR data_array.data0\[12\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_138_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11818_ clknet_leaf_126_clk _00626_ VGND VGND VPWR VPWR data_array.data0\[7\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_12798_ clknet_leaf_135_clk _01492_ VGND VGND VPWR VPWR tag_array.tag1\[10\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_61_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11749_ clknet_leaf_64_clk _00557_ VGND VGND VPWR VPWR data_array.data0\[8\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_159_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14468_ clknet_leaf_211_clk _03091_ VGND VGND VPWR VPWR data_array.data1\[7\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
X_13419_ clknet_leaf_240_clk _02049_ VGND VGND VPWR VPWR data_array.data1\[8\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_155_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14399_ clknet_leaf_40_clk _03022_ VGND VGND VPWR VPWR data_array.data1\[10\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_154_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08960_ net927 net2903 net426 VGND VGND VPWR VPWR _00716_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_5_clk clknet_5_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07911_ net1631 _05103_ _05107_ net1205 VGND VGND VPWR VPWR _05110_ sky130_fd_sc_hd__a22o_1
Xhold2506 tag_array.tag0\[11\]\[5\] VGND VGND VPWR VPWR net4157 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2517 data_array.data1\[9\]\[48\] VGND VGND VPWR VPWR net4168 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08891_ net940 net4113 net440 VGND VGND VPWR VPWR _00648_ sky130_fd_sc_hd__mux2_1
Xhold2528 tag_array.tag0\[2\]\[7\] VGND VGND VPWR VPWR net4179 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_16_Left_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2539 data_array.data1\[9\]\[50\] VGND VGND VPWR VPWR net4190 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_64_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1805 data_array.data1\[10\]\[23\] VGND VGND VPWR VPWR net3456 sky130_fd_sc_hd__dlygate4sd3_1
X_07842_ data_array.data1\[12\]\[36\] net1416 net1322 data_array.data1\[15\]\[36\]
+ _05046_ VGND VGND VPWR VPWR _05047_ sky130_fd_sc_hd__a221o_1
Xhold1816 data_array.data1\[2\]\[35\] VGND VGND VPWR VPWR net3467 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1827 data_array.data1\[5\]\[28\] VGND VGND VPWR VPWR net3478 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1838 data_array.data0\[5\]\[14\] VGND VGND VPWR VPWR net3489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1849 tag_array.tag1\[7\]\[24\] VGND VGND VPWR VPWR net3500 sky130_fd_sc_hd__dlygate4sd3_1
X_07773_ data_array.data1\[5\]\[30\] net1583 net1487 data_array.data1\[6\]\[30\] VGND
+ VGND VPWR VPWR _04984_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_179_3800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclone8 net853 VGND VGND VPWR VPWR net1659 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09512_ net781 net3152 net621 VGND VGND VPWR VPWR _01265_ sky130_fd_sc_hd__mux2_1
X_06724_ net1185 _04025_ _04029_ net1233 VGND VGND VPWR VPWR _04031_ sky130_fd_sc_hd__a22o_1
XFILLER_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09443_ net892 net3428 net579 VGND VGND VPWR VPWR _01196_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_175_3719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06655_ tag_array.tag1\[1\]\[17\] net1607 net1511 tag_array.tag1\[2\]\[17\] VGND
+ VGND VPWR VPWR _03968_ sky130_fd_sc_hd__a22o_1
XFILLER_25_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09374_ net904 net4431 net402 VGND VGND VPWR VPWR _01127_ sky130_fd_sc_hd__mux2_1
X_06586_ tag_array.tag1\[4\]\[11\] net1388 net1294 tag_array.tag1\[7\]\[11\] _03904_
+ VGND VGND VPWR VPWR _03905_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_25_Left_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08325_ net107 net42 net1639 VGND VGND VPWR VPWR _05453_ sky130_fd_sc_hd__mux2_1
XFILLER_21_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08256_ net711 net3584 net796 VGND VGND VPWR VPWR _00216_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_468 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07207_ net1631 _04463_ _04467_ net1205 VGND VGND VPWR VPWR _04470_ sky130_fd_sc_hd__a22o_1
X_08187_ net1649 net1159 fsm.lru_out VGND VGND VPWR VPWR _05357_ sky130_fd_sc_hd__and3_1
XFILLER_165_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07138_ data_array.data0\[12\]\[36\] net1413 net1319 data_array.data0\[15\]\[36\]
+ _04406_ VGND VGND VPWR VPWR _04407_ sky130_fd_sc_hd__a221o_1
XFILLER_152_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07069_ data_array.data0\[5\]\[30\] net1582 net1486 data_array.data0\[6\]\[30\] VGND
+ VGND VPWR VPWR _04344_ sky130_fd_sc_hd__a22o_1
XFILLER_121_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput260 net260 VGND VGND VPWR VPWR mem_addr[8] sky130_fd_sc_hd__buf_2
XFILLER_0_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput271 net271 VGND VGND VPWR VPWR mem_wdata[17] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput282 net282 VGND VGND VPWR VPWR mem_wdata[27] sky130_fd_sc_hd__buf_2
Xoutput293 net293 VGND VGND VPWR VPWR mem_wdata[37] sky130_fd_sc_hd__buf_2
XFILLER_59_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10080_ net705 net2579 net601 VGND VGND VPWR VPWR _01829_ sky130_fd_sc_hd__mux2_1
XFILLER_181_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13770_ clknet_leaf_253_clk _02399_ VGND VGND VPWR VPWR data_array.data1\[2\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_43_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10982_ net2137 net1072 net341 VGND VGND VPWR VPWR _02726_ sky130_fd_sc_hd__mux2_1
XFILLER_43_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12721_ clknet_leaf_169_clk _01415_ VGND VGND VPWR VPWR tag_array.tag0\[7\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12652_ clknet_leaf_10_clk _01346_ VGND VGND VPWR VPWR data_array.data0\[15\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
X_11603_ clknet_leaf_95_clk _00411_ VGND VGND VPWR VPWR tag_array.tag1\[4\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_12583_ clknet_leaf_162_clk _01277_ VGND VGND VPWR VPWR tag_array.tag0\[10\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_169_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14322_ clknet_leaf_88_clk _02951_ VGND VGND VPWR VPWR data_array.data1\[11\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_157_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11534_ clknet_leaf_97_clk _00342_ VGND VGND VPWR VPWR tag_array.tag1\[6\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_184_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_150_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14253_ clknet_leaf_217_clk _02882_ VGND VGND VPWR VPWR data_array.data1\[12\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_20 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11465_ clknet_leaf_221_clk _00275_ VGND VGND VPWR VPWR data_array.data0\[0\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
X_13204_ clknet_leaf_256_clk _00099_ VGND VGND VPWR VPWR data_array.rdata1\[41\] sky130_fd_sc_hd__dfxtp_1
X_10416_ net2252 net990 net668 VGND VGND VPWR VPWR _02162_ sky130_fd_sc_hd__mux2_1
X_14184_ clknet_leaf_258_clk _02813_ VGND VGND VPWR VPWR data_array.data0\[2\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_74_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11396_ clknet_leaf_103_clk _00206_ VGND VGND VPWR VPWR tag_array.tag1\[7\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_152_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13135_ clknet_leaf_190_clk _01829_ VGND VGND VPWR VPWR tag_array.tag0\[3\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_10347_ net712 net4153 net591 VGND VGND VPWR VPWR _02094_ sky130_fd_sc_hd__mux2_1
XFILLER_3_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13066_ clknet_leaf_255_clk _01760_ VGND VGND VPWR VPWR data_array.data1\[13\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_10278_ net2183 net1050 net640 VGND VGND VPWR VPWR _02025_ sky130_fd_sc_hd__mux2_1
Xfanout1430 net1434 VGND VGND VPWR VPWR net1430 sky130_fd_sc_hd__clkbuf_4
X_12017_ clknet_leaf_239_clk _00825_ VGND VGND VPWR VPWR data_array.data0\[6\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout1441 net1443 VGND VGND VPWR VPWR net1441 sky130_fd_sc_hd__clkbuf_4
XFILLER_79_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1452 net1453 VGND VGND VPWR VPWR net1452 sky130_fd_sc_hd__clkbuf_4
XFILLER_39_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1463 net1464 VGND VGND VPWR VPWR net1463 sky130_fd_sc_hd__clkbuf_4
Xfanout1474 net1477 VGND VGND VPWR VPWR net1474 sky130_fd_sc_hd__clkbuf_4
Xfanout1485 net1486 VGND VGND VPWR VPWR net1485 sky130_fd_sc_hd__clkbuf_4
Xfanout1496 net1498 VGND VGND VPWR VPWR net1496 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13968_ clknet_leaf_28_clk _02597_ VGND VGND VPWR VPWR data_array.data1\[5\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1024 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12919_ clknet_leaf_176_clk _01613_ VGND VGND VPWR VPWR data_array.data0\[13\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13899_ clknet_leaf_28_clk _02528_ VGND VGND VPWR VPWR data_array.data1\[4\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_06440_ tag_array.tag0\[9\]\[23\] net1607 net1511 tag_array.tag0\[10\]\[23\] VGND
+ VGND VPWR VPWR _03772_ sky130_fd_sc_hd__a22o_1
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06371_ net1634 _03703_ _03707_ net1208 VGND VGND VPWR VPWR _03710_ sky130_fd_sc_hd__a22o_1
XFILLER_175_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_170_3627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08110_ net1183 _05285_ _05289_ net1233 VGND VGND VPWR VPWR _05291_ sky130_fd_sc_hd__a22o_1
XFILLER_148_958 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09090_ net927 net4588 net410 VGND VGND VPWR VPWR _00844_ sky130_fd_sc_hd__mux2_1
XFILLER_30_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08041_ data_array.data1\[5\]\[54\] net1544 net1448 data_array.data1\[6\]\[54\] VGND
+ VGND VPWR VPWR _05228_ sky130_fd_sc_hd__a22o_1
XFILLER_31_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold902 data_array.data0\[5\]\[57\] VGND VGND VPWR VPWR net2553 sky130_fd_sc_hd__dlygate4sd3_1
Xhold913 tag_array.tag0\[15\]\[11\] VGND VGND VPWR VPWR net2564 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_31_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold924 data_array.data1\[13\]\[36\] VGND VGND VPWR VPWR net2575 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold935 data_array.data0\[13\]\[12\] VGND VGND VPWR VPWR net2586 sky130_fd_sc_hd__dlygate4sd3_1
Xhold946 tag_array.tag0\[9\]\[21\] VGND VGND VPWR VPWR net2597 sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 data_array.data1\[9\]\[3\] VGND VGND VPWR VPWR net2608 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold968 data_array.data1\[12\]\[13\] VGND VGND VPWR VPWR net2619 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_354 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09992_ net860 net2612 net377 VGND VGND VPWR VPWR _01741_ sky130_fd_sc_hd__mux2_1
XFILLER_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold979 data_array.data1\[1\]\[1\] VGND VGND VPWR VPWR net2630 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_168_3589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08943_ net992 net3728 net430 VGND VGND VPWR VPWR _00699_ sky130_fd_sc_hd__mux2_1
Xhold2303 tag_array.tag1\[15\]\[12\] VGND VGND VPWR VPWR net3954 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2314 tag_array.tag1\[6\]\[10\] VGND VGND VPWR VPWR net3965 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2325 data_array.data0\[7\]\[13\] VGND VGND VPWR VPWR net3976 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_4_15_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_15_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_32_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2336 data_array.data0\[14\]\[34\] VGND VGND VPWR VPWR net3987 sky130_fd_sc_hd__dlygate4sd3_1
X_08874_ net1009 net4214 net434 VGND VGND VPWR VPWR _00631_ sky130_fd_sc_hd__mux2_1
XFILLER_57_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1602 tag_array.tag0\[6\]\[8\] VGND VGND VPWR VPWR net3253 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2347 tag_array.tag0\[4\]\[0\] VGND VGND VPWR VPWR net3998 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1613 data_array.data0\[11\]\[40\] VGND VGND VPWR VPWR net3264 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2358 data_array.data1\[7\]\[6\] VGND VGND VPWR VPWR net4009 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1624 data_array.data1\[12\]\[1\] VGND VGND VPWR VPWR net3275 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2369 tag_array.tag1\[14\]\[2\] VGND VGND VPWR VPWR net4020 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1635 tag_array.tag1\[2\]\[20\] VGND VGND VPWR VPWR net3286 sky130_fd_sc_hd__dlygate4sd3_1
X_07825_ _05030_ _05031_ VGND VGND VPWR VPWR _00091_ sky130_fd_sc_hd__or2_1
XFILLER_57_647 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1646 data_array.data0\[12\]\[33\] VGND VGND VPWR VPWR net3297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1657 data_array.data1\[2\]\[6\] VGND VGND VPWR VPWR net3308 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1668 tag_array.tag1\[14\]\[21\] VGND VGND VPWR VPWR net3319 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1679 data_array.data0\[14\]\[11\] VGND VGND VPWR VPWR net3330 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07756_ data_array.data1\[0\]\[28\] net1349 net1255 data_array.data1\[3\]\[28\] _04968_
+ VGND VGND VPWR VPWR _04969_ sky130_fd_sc_hd__a221o_1
X_06707_ tag_array.tag1\[0\]\[22\] net1362 net1268 tag_array.tag1\[3\]\[22\] _04014_
+ VGND VGND VPWR VPWR _04015_ sky130_fd_sc_hd__a221o_1
X_07687_ data_array.data1\[13\]\[22\] net1539 net1443 data_array.data1\[14\]\[22\]
+ VGND VGND VPWR VPWR _04906_ sky130_fd_sc_hd__a22o_1
X_09426_ net962 net3882 net582 VGND VGND VPWR VPWR _01179_ sky130_fd_sc_hd__mux2_1
X_06638_ tag_array.tag1\[13\]\[16\] net1609 net1513 tag_array.tag1\[14\]\[16\] VGND
+ VGND VPWR VPWR _03952_ sky130_fd_sc_hd__a22o_1
XFILLER_53_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09357_ net973 net3987 net402 VGND VGND VPWR VPWR _01110_ sky130_fd_sc_hd__mux2_1
X_06569_ net1636 _03883_ _03887_ net1210 VGND VGND VPWR VPWR _03890_ sky130_fd_sc_hd__a22o_1
XFILLER_138_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08308_ net1128 _05441_ VGND VGND VPWR VPWR _05442_ sky130_fd_sc_hd__and2_1
X_09288_ net728 net3307 net564 VGND VGND VPWR VPWR _01042_ sky130_fd_sc_hd__mux2_1
XFILLER_138_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08239_ net1651 net1161 net15 VGND VGND VPWR VPWR _05394_ sky130_fd_sc_hd__and3_1
XFILLER_119_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11250_ net1031 net3346 net683 VGND VGND VPWR VPWR _02993_ sky130_fd_sc_hd__mux2_1
XFILLER_153_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10201_ net1002 net4404 net357 VGND VGND VPWR VPWR _01948_ sky130_fd_sc_hd__mux2_1
X_11181_ net1050 net3358 net656 VGND VGND VPWR VPWR _02924_ sky130_fd_sc_hd__mux2_1
XFILLER_106_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10132_ net1018 net3682 net364 VGND VGND VPWR VPWR _01880_ sky130_fd_sc_hd__mux2_1
XFILLER_121_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10063_ net771 net4038 net600 VGND VGND VPWR VPWR _01812_ sky130_fd_sc_hd__mux2_1
XFILLER_76_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2870 data_array.data1\[13\]\[35\] VGND VGND VPWR VPWR net4521 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2881 data_array.data0\[14\]\[24\] VGND VGND VPWR VPWR net4532 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2892 data_array.data1\[14\]\[38\] VGND VGND VPWR VPWR net4543 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13822_ clknet_leaf_215_clk _02451_ VGND VGND VPWR VPWR data_array.data1\[2\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13753_ clknet_leaf_55_clk _02382_ VGND VGND VPWR VPWR data_array.data1\[1\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
X_10965_ net883 net2754 net526 VGND VGND VPWR VPWR _02710_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12704_ clknet_leaf_185_clk _01398_ VGND VGND VPWR VPWR tag_array.tag0\[8\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_104_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13684_ clknet_leaf_82_clk _02313_ VGND VGND VPWR VPWR data_array.data1\[15\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
X_10896_ net900 net2697 net516 VGND VGND VPWR VPWR _02641_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_84_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12635_ clknet_leaf_249_clk _01329_ VGND VGND VPWR VPWR data_array.data0\[15\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12566_ clknet_leaf_143_clk _01260_ VGND VGND VPWR VPWR tag_array.tag0\[11\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_79_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11517_ clknet_leaf_135_clk _00325_ VGND VGND VPWR VPWR tag_array.tag1\[9\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_14305_ clknet_leaf_268_clk _02934_ VGND VGND VPWR VPWR data_array.data1\[11\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12497_ clknet_leaf_40_clk _01191_ VGND VGND VPWR VPWR data_array.data1\[9\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
X_14236_ clknet_leaf_130_clk _02865_ VGND VGND VPWR VPWR data_array.data1\[12\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold209 data_array.data0\[8\]\[43\] VGND VGND VPWR VPWR net1860 sky130_fd_sc_hd__dlygate4sd3_1
X_11448_ clknet_leaf_217_clk _00258_ VGND VGND VPWR VPWR data_array.data0\[0\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14167_ clknet_leaf_63_clk _02796_ VGND VGND VPWR VPWR data_array.data0\[2\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_11379_ net819 net3373 _05578_ VGND VGND VPWR VPWR _03122_ sky130_fd_sc_hd__mux2_1
XFILLER_140_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13118_ clknet_leaf_141_clk _01812_ VGND VGND VPWR VPWR tag_array.tag0\[3\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_14098_ clknet_leaf_112_clk _02727_ VGND VGND VPWR VPWR data_array.data0\[1\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_05940_ data_array.rdata1\[36\] net1657 net843 VGND VGND VPWR VPWR _03421_ sky130_fd_sc_hd__a21o_1
XFILLER_39_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13049_ clknet_leaf_226_clk _01743_ VGND VGND VPWR VPWR data_array.data1\[13\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1260 net1261 VGND VGND VPWR VPWR net1260 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_163_3486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1271 net1273 VGND VGND VPWR VPWR net1271 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_163_3497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05871_ data_array.rdata1\[13\] net831 net840 VGND VGND VPWR VPWR _03375_ sky130_fd_sc_hd__a21o_1
XFILLER_38_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1282 _03515_ VGND VGND VPWR VPWR net1282 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_1_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1293 net1294 VGND VGND VPWR VPWR net1293 sky130_fd_sc_hd__clkbuf_4
X_07610_ data_array.data1\[13\]\[15\] net1581 net1485 data_array.data1\[14\]\[15\]
+ VGND VGND VPWR VPWR _04836_ sky130_fd_sc_hd__a22o_1
XFILLER_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08590_ net764 net4516 net536 VGND VGND VPWR VPWR _00349_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_124_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07541_ data_array.data1\[8\]\[9\] net1391 net1297 data_array.data1\[11\]\[9\] _04772_
+ VGND VGND VPWR VPWR _04773_ sky130_fd_sc_hd__a221o_1
XFILLER_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07472_ net1166 _04705_ _04709_ net1214 VGND VGND VPWR VPWR _04711_ sky130_fd_sc_hd__a22o_1
X_09211_ net736 net3177 net630 VGND VGND VPWR VPWR _00965_ sky130_fd_sc_hd__mux2_1
XFILLER_179_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06423_ tag_array.tag0\[8\]\[21\] net1408 net1314 tag_array.tag0\[11\]\[21\] _03756_
+ VGND VGND VPWR VPWR _03757_ sky130_fd_sc_hd__a221o_1
XFILLER_50_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09142_ net974 net3972 net568 VGND VGND VPWR VPWR _00896_ sky130_fd_sc_hd__mux2_1
X_06354_ tag_array.tag0\[1\]\[15\] net1593 net1497 tag_array.tag0\[2\]\[15\] VGND
+ VGND VPWR VPWR _03694_ sky130_fd_sc_hd__a22o_1
X_09073_ net992 net4488 net414 VGND VGND VPWR VPWR _00827_ sky130_fd_sc_hd__mux2_1
X_06285_ _03630_ _03631_ VGND VGND VPWR VPWR _00154_ sky130_fd_sc_hd__or2_1
X_08024_ data_array.data1\[9\]\[53\] net1523 net1427 data_array.data1\[10\]\[53\]
+ VGND VGND VPWR VPWR _05212_ sky130_fd_sc_hd__a22o_1
XFILLER_135_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold710 data_array.data0\[12\]\[62\] VGND VGND VPWR VPWR net2361 sky130_fd_sc_hd__dlygate4sd3_1
Xhold721 data_array.data1\[0\]\[21\] VGND VGND VPWR VPWR net2372 sky130_fd_sc_hd__dlygate4sd3_1
Xhold732 tag_array.tag1\[15\]\[15\] VGND VGND VPWR VPWR net2383 sky130_fd_sc_hd__dlygate4sd3_1
Xhold743 data_array.data0\[12\]\[5\] VGND VGND VPWR VPWR net2394 sky130_fd_sc_hd__dlygate4sd3_1
Xhold754 data_array.data0\[12\]\[31\] VGND VGND VPWR VPWR net2405 sky130_fd_sc_hd__dlygate4sd3_1
Xhold765 tag_array.tag1\[10\]\[5\] VGND VGND VPWR VPWR net2416 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold776 data_array.data1\[15\]\[34\] VGND VGND VPWR VPWR net2427 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_536 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold787 tag_array.tag0\[15\]\[8\] VGND VGND VPWR VPWR net2438 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold798 data_array.data0\[6\]\[6\] VGND VGND VPWR VPWR net2449 sky130_fd_sc_hd__dlygate4sd3_1
X_09975_ net928 net4134 net371 VGND VGND VPWR VPWR _01724_ sky130_fd_sc_hd__mux2_1
XFILLER_89_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2100 data_array.data1\[7\]\[55\] VGND VGND VPWR VPWR net3751 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2111 lru_array.lru_mem\[11\] VGND VGND VPWR VPWR net3762 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2122 data_array.data1\[13\]\[63\] VGND VGND VPWR VPWR net3773 sky130_fd_sc_hd__dlygate4sd3_1
X_08926_ net1060 net3282 net432 VGND VGND VPWR VPWR _00682_ sky130_fd_sc_hd__mux2_1
XFILLER_58_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2133 tag_array.tag0\[9\]\[5\] VGND VGND VPWR VPWR net3784 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2144 data_array.data1\[3\]\[58\] VGND VGND VPWR VPWR net3795 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1410 tag_array.tag0\[11\]\[3\] VGND VGND VPWR VPWR net3061 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2155 lru_array.lru_mem\[13\] VGND VGND VPWR VPWR net3806 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1421 data_array.data0\[12\]\[41\] VGND VGND VPWR VPWR net3072 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2166 data_array.data1\[5\]\[13\] VGND VGND VPWR VPWR net3817 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2177 tag_array.tag0\[1\]\[3\] VGND VGND VPWR VPWR net3828 sky130_fd_sc_hd__dlygate4sd3_1
X_08857_ net1076 net3468 net434 VGND VGND VPWR VPWR _00614_ sky130_fd_sc_hd__mux2_1
Xhold1432 tag_array.tag0\[2\]\[5\] VGND VGND VPWR VPWR net3083 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1443 data_array.data1\[10\]\[25\] VGND VGND VPWR VPWR net3094 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2188 tag_array.tag0\[3\]\[3\] VGND VGND VPWR VPWR net3839 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2199 data_array.data1\[12\]\[36\] VGND VGND VPWR VPWR net3850 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1454 data_array.data0\[12\]\[0\] VGND VGND VPWR VPWR net3105 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1465 tag_array.tag0\[13\]\[3\] VGND VGND VPWR VPWR net3116 sky130_fd_sc_hd__dlygate4sd3_1
X_07808_ data_array.data1\[9\]\[33\] net1588 net1492 data_array.data1\[10\]\[33\]
+ VGND VGND VPWR VPWR _05016_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_220_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_220_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold1476 data_array.data0\[15\]\[26\] VGND VGND VPWR VPWR net3127 sky130_fd_sc_hd__dlygate4sd3_1
X_08788_ net3214 net1093 net446 VGND VGND VPWR VPWR _00546_ sky130_fd_sc_hd__mux2_1
Xhold1487 tag_array.tag0\[12\]\[13\] VGND VGND VPWR VPWR net3138 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1498 tag_array.tag0\[2\]\[15\] VGND VGND VPWR VPWR net3149 sky130_fd_sc_hd__dlygate4sd3_1
X_07739_ data_array.data1\[8\]\[27\] net1358 net1264 data_array.data1\[11\]\[27\]
+ _04952_ VGND VGND VPWR VPWR _04953_ sky130_fd_sc_hd__a221o_1
XFILLER_77_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10750_ net974 net3067 net492 VGND VGND VPWR VPWR _02495_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_9_Left_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09409_ net1031 net3124 net588 VGND VGND VPWR VPWR _01162_ sky130_fd_sc_hd__mux2_1
XFILLER_52_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10681_ net3334 net995 net483 VGND VGND VPWR VPWR _02426_ sky130_fd_sc_hd__mux2_1
XFILLER_139_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12420_ clknet_leaf_73_clk _01114_ VGND VGND VPWR VPWR data_array.data0\[14\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_62_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12351_ clknet_leaf_77_clk _00026_ VGND VGND VPWR VPWR data_array.rdata0\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11302_ net1086 net4009 net795 VGND VGND VPWR VPWR _03045_ sky130_fd_sc_hd__mux2_1
XFILLER_14_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12282_ clknet_leaf_231_clk _01040_ VGND VGND VPWR VPWR tag_array.tag1\[13\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14021_ clknet_leaf_211_clk _02650_ VGND VGND VPWR VPWR data_array.data1\[5\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_181_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11233_ net1099 net3715 net675 VGND VGND VPWR VPWR _02976_ sky130_fd_sc_hd__mux2_1
XFILLER_84_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11164_ net863 net3578 net551 VGND VGND VPWR VPWR _02907_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10115_ net1084 net3496 net362 VGND VGND VPWR VPWR _01863_ sky130_fd_sc_hd__mux2_1
XFILLER_49_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_817 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11095_ net3662 net880 net332 VGND VGND VPWR VPWR _02838_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_145_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10046_ net901 net2530 net558 VGND VGND VPWR VPWR _01795_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_69_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold70 tag_array.valid0\[9\] VGND VGND VPWR VPWR net1721 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_211_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_211_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold81 tag_array.tag1\[1\]\[18\] VGND VGND VPWR VPWR net1732 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 data_array.data1\[2\]\[15\] VGND VGND VPWR VPWR net1743 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_36_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_141_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13805_ clknet_leaf_214_clk _02434_ VGND VGND VPWR VPWR data_array.data1\[2\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
X_11997_ clknet_leaf_104_clk _00805_ VGND VGND VPWR VPWR data_array.data0\[6\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10948_ net950 net2753 net535 VGND VGND VPWR VPWR _02693_ sky130_fd_sc_hd__mux2_1
XFILLER_17_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13736_ clknet_leaf_257_clk _02365_ VGND VGND VPWR VPWR data_array.data1\[1\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_82_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10879_ net968 net3037 net515 VGND VGND VPWR VPWR _02624_ sky130_fd_sc_hd__mux2_1
X_13667_ clknet_leaf_221_clk _02296_ VGND VGND VPWR VPWR data_array.data1\[15\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_12618_ clknet_leaf_230_clk _01312_ VGND VGND VPWR VPWR data_array.data0\[15\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_13598_ clknet_leaf_192_clk _02227_ VGND VGND VPWR VPWR data_array.data0\[9\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_157_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12549_ clknet_leaf_179_clk _01243_ VGND VGND VPWR VPWR tag_array.tag0\[11\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_1 _00002_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06070_ fsm.tag_out0\[17\] net1121 _03498_ VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__a21o_1
XFILLER_133_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14219_ clknet_leaf_35_clk _02848_ VGND VGND VPWR VPWR data_array.data1\[12\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_165_3526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_3537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout508 net512 VGND VGND VPWR VPWR net508 sky130_fd_sc_hd__clkbuf_8
Xfanout519 net522 VGND VGND VPWR VPWR net519 sky130_fd_sc_hd__clkbuf_8
X_09760_ net2270 net746 net670 VGND VGND VPWR VPWR _01512_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_182_3851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06972_ data_array.data0\[13\]\[21\] net1556 net1460 data_array.data0\[14\]\[21\]
+ VGND VGND VPWR VPWR _04256_ sky130_fd_sc_hd__a22o_1
XFILLER_140_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_182_3862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08711_ net2160 net778 net470 VGND VGND VPWR VPWR _00470_ sky130_fd_sc_hd__mux2_1
X_05923_ net122 net1155 _03408_ _03409_ VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__a22o_1
XFILLER_39_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09691_ net722 net4344 net606 VGND VGND VPWR VPWR _01443_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_202_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_202_clk
+ sky130_fd_sc_hd__clkbuf_8
Xfanout1090 net1091 VGND VGND VPWR VPWR net1090 sky130_fd_sc_hd__clkbuf_2
XFILLER_27_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08642_ net4461 net756 net510 VGND VGND VPWR VPWR _00401_ sky130_fd_sc_hd__mux2_1
X_05854_ net160 net1157 _03362_ _03363_ VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__a22o_1
XFILLER_94_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08573_ net811 _05583_ net1696 VGND VGND VPWR VPWR _00337_ sky130_fd_sc_hd__a21o_1
X_05785_ net15 _03141_ _03257_ _03300_ _03301_ VGND VGND VPWR VPWR _03302_ sky130_fd_sc_hd__a2111o_1
XFILLER_23_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07524_ data_array.data1\[5\]\[7\] net1589 net1493 data_array.data1\[6\]\[7\] VGND
+ VGND VPWR VPWR _04758_ sky130_fd_sc_hd__a22o_1
X_07455_ data_array.data1\[0\]\[1\] net1330 net1236 data_array.data1\[3\]\[1\] _04694_
+ VGND VGND VPWR VPWR _04695_ sky130_fd_sc_hd__a221o_1
X_06406_ _03740_ _03741_ VGND VGND VPWR VPWR _00141_ sky130_fd_sc_hd__or2_1
XFILLER_50_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07386_ data_array.data0\[9\]\[59\] net1570 net1474 data_array.data0\[10\]\[59\]
+ VGND VGND VPWR VPWR _04632_ sky130_fd_sc_hd__a22o_1
XFILLER_148_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09125_ net1041 net2228 net567 VGND VGND VPWR VPWR _00879_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_269_clk clknet_5_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_269_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_157_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06337_ tag_array.tag0\[4\]\[13\] net1417 net1323 tag_array.tag0\[7\]\[13\] _03678_
+ VGND VGND VPWR VPWR _03679_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_40_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09056_ net1060 net3410 net416 VGND VGND VPWR VPWR _00810_ sky130_fd_sc_hd__mux2_1
X_06268_ tag_array.tag0\[13\]\[7\] net1598 net1502 tag_array.tag0\[14\]\[7\] VGND
+ VGND VPWR VPWR _03616_ sky130_fd_sc_hd__a22o_1
XFILLER_135_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08007_ data_array.data1\[8\]\[51\] net1334 net1240 data_array.data1\[11\]\[51\]
+ _05196_ VGND VGND VPWR VPWR _05197_ sky130_fd_sc_hd__a221o_1
XFILLER_135_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold540 data_array.data1\[4\]\[27\] VGND VGND VPWR VPWR net2191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold551 data_array.data0\[14\]\[40\] VGND VGND VPWR VPWR net2202 sky130_fd_sc_hd__dlygate4sd3_1
X_06199_ tag_array.tag0\[8\]\[1\] net1402 net1308 tag_array.tag0\[11\]\[1\] _03552_
+ VGND VGND VPWR VPWR _03553_ sky130_fd_sc_hd__a221o_1
XFILLER_117_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold562 data_array.data1\[4\]\[46\] VGND VGND VPWR VPWR net2213 sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 data_array.data1\[0\]\[35\] VGND VGND VPWR VPWR net2224 sky130_fd_sc_hd__dlygate4sd3_1
Xhold584 data_array.data1\[2\]\[51\] VGND VGND VPWR VPWR net2235 sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 tag_array.tag1\[0\]\[3\] VGND VGND VPWR VPWR net2246 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09958_ net996 net3787 net371 VGND VGND VPWR VPWR _01707_ sky130_fd_sc_hd__mux2_1
X_08909_ net868 net2639 net440 VGND VGND VPWR VPWR _00666_ sky130_fd_sc_hd__mux2_1
XFILLER_106_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09889_ net913 net2165 net383 VGND VGND VPWR VPWR _01639_ sky130_fd_sc_hd__mux2_1
Xhold1240 data_array.data1\[2\]\[48\] VGND VGND VPWR VPWR net2891 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1251 data_array.data1\[5\]\[30\] VGND VGND VPWR VPWR net2902 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_872 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1262 tag_array.tag1\[8\]\[5\] VGND VGND VPWR VPWR net2913 sky130_fd_sc_hd__dlygate4sd3_1
X_11920_ clknet_leaf_208_clk _00728_ VGND VGND VPWR VPWR data_array.data0\[5\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_131_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1273 data_array.data0\[4\]\[38\] VGND VGND VPWR VPWR net2924 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_174_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1284 tag_array.tag0\[6\]\[15\] VGND VGND VPWR VPWR net2935 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1295 data_array.data0\[12\]\[22\] VGND VGND VPWR VPWR net2946 sky130_fd_sc_hd__dlygate4sd3_1
X_11851_ clknet_leaf_2_clk _00659_ VGND VGND VPWR VPWR data_array.data0\[7\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10802_ net1901 net1021 net503 VGND VGND VPWR VPWR _02547_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11782_ clknet_leaf_90_clk _00590_ VGND VGND VPWR VPWR data_array.data0\[8\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
X_10733_ net1040 net4478 net490 VGND VGND VPWR VPWR _02478_ sky130_fd_sc_hd__mux2_1
X_13521_ clknet_leaf_18_clk _02150_ VGND VGND VPWR VPWR data_array.data1\[0\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_24_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13452_ clknet_leaf_144_clk _02082_ VGND VGND VPWR VPWR tag_array.tag0\[1\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_10664_ net2781 net1062 net484 VGND VGND VPWR VPWR _02409_ sky130_fd_sc_hd__mux2_1
XFILLER_90_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12403_ clknet_leaf_226_clk _01097_ VGND VGND VPWR VPWR data_array.data0\[14\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_166_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13383_ clknet_leaf_28_clk _02013_ VGND VGND VPWR VPWR data_array.data1\[8\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_167_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10595_ net1804 net1083 net473 VGND VGND VPWR VPWR _02340_ sky130_fd_sc_hd__mux2_1
X_12334_ clknet_leaf_212_clk _00007_ VGND VGND VPWR VPWR data_array.rdata0\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_115_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12265_ clknet_leaf_196_clk _01023_ VGND VGND VPWR VPWR tag_array.tag1\[14\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_587 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_128_Right_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14004_ clknet_leaf_84_clk _02633_ VGND VGND VPWR VPWR data_array.data1\[5\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
X_11216_ net910 net2509 net649 VGND VGND VPWR VPWR _02959_ sky130_fd_sc_hd__mux2_1
XFILLER_122_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12196_ clknet_leaf_182_clk _00149_ VGND VGND VPWR VPWR fsm.tag_out0\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_150_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11147_ net931 net2745 net543 VGND VGND VPWR VPWR _02890_ sky130_fd_sc_hd__mux2_1
XFILLER_110_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_143_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11078_ net1755 net948 net335 VGND VGND VPWR VPWR _02821_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_160_3434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput160 mem_rdata[7] VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_160_3445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10029_ net969 net4521 net554 VGND VGND VPWR VPWR _01778_ sky130_fd_sc_hd__mux2_1
XFILLER_64_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13719_ clknet_leaf_64_clk _02348_ VGND VGND VPWR VPWR data_array.data1\[1\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_158_3396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07240_ net1192 _04493_ _04497_ net1618 VGND VGND VPWR VPWR _04500_ sky130_fd_sc_hd__a22o_1
XFILLER_32_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07171_ data_array.data0\[12\]\[39\] net1349 net1255 data_array.data0\[15\]\[39\]
+ _04436_ VGND VGND VPWR VPWR _04437_ sky130_fd_sc_hd__a221o_1
XFILLER_157_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06122_ data_array.rdata0\[37\] net1136 net1117 data_array.rdata1\[37\] VGND VGND
+ VPWR VPWR net293 sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_136_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06053_ net1163 net8 fsm.tag_out1\[9\] net1132 VGND VGND VPWR VPWR _03490_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_184_3902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_184_3913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_1054 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09812_ net961 net3339 net388 VGND VGND VPWR VPWR _01563_ sky130_fd_sc_hd__mux2_1
XFILLER_86_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout338 net339 VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__buf_4
XFILLER_87_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout349 net350 VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__buf_4
XFILLER_115_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06955_ net1180 _04235_ _04239_ net1226 VGND VGND VPWR VPWR _04241_ sky130_fd_sc_hd__a22o_1
X_09743_ net715 net4266 net680 VGND VGND VPWR VPWR _01495_ sky130_fd_sc_hd__mux2_1
X_05906_ data_array.rdata0\[25\] net846 net1142 VGND VGND VPWR VPWR _03398_ sky130_fd_sc_hd__o21a_1
X_09674_ net793 net3160 net606 VGND VGND VPWR VPWR _01426_ sky130_fd_sc_hd__mux2_1
X_06886_ data_array.data0\[5\]\[13\] net1549 net1453 data_array.data0\[6\]\[13\] VGND
+ VGND VPWR VPWR _04178_ sky130_fd_sc_hd__a22o_1
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08625_ net724 net3701 net523 VGND VGND VPWR VPWR _00384_ sky130_fd_sc_hd__mux2_1
XFILLER_54_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05837_ data_array.rdata0\[2\] net848 net1142 VGND VGND VPWR VPWR _03352_ sky130_fd_sc_hd__o21a_1
XFILLER_70_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08556_ net731 net4535 net585 VGND VGND VPWR VPWR _00324_ sky130_fd_sc_hd__mux2_1
X_05768_ _03241_ _03255_ _03268_ _03284_ VGND VGND VPWR VPWR _03285_ sky130_fd_sc_hd__or4_1
X_07507_ data_array.data1\[9\]\[6\] net1519 net1423 data_array.data1\[10\]\[6\] VGND
+ VGND VPWR VPWR _04742_ sky130_fd_sc_hd__a22o_1
XFILLER_168_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08487_ _03514_ _03523_ VGND VGND VPWR VPWR _05561_ sky130_fd_sc_hd__nor2_1
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05699_ _03142_ fsm.tag_out0\[18\] _03172_ _03178_ net1654 VGND VGND VPWR VPWR _03216_
+ sky130_fd_sc_hd__a2111o_1
XFILLER_168_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07438_ net1198 _04673_ _04677_ net1624 VGND VGND VPWR VPWR _04680_ sky130_fd_sc_hd__a22o_1
XFILLER_10_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07369_ data_array.data0\[8\]\[57\] net1347 net1253 data_array.data0\[11\]\[57\]
+ _04616_ VGND VGND VPWR VPWR _04617_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_99_Left_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09108_ net1111 net2864 net571 VGND VGND VPWR VPWR _00862_ sky130_fd_sc_hd__mux2_1
XFILLER_109_758 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10380_ net353 net3084 net557 VGND VGND VPWR VPWR _02126_ sky130_fd_sc_hd__mux2_1
XFILLER_108_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09039_ net1990 net868 net424 VGND VGND VPWR VPWR _00794_ sky130_fd_sc_hd__mux2_1
XFILLER_184_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12050_ clknet_leaf_110_clk _00858_ VGND VGND VPWR VPWR data_array.data0\[6\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold370 data_array.data1\[8\]\[25\] VGND VGND VPWR VPWR net2021 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold381 data_array.data1\[4\]\[57\] VGND VGND VPWR VPWR net2032 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold392 data_array.data0\[0\]\[2\] VGND VGND VPWR VPWR net2043 sky130_fd_sc_hd__dlygate4sd3_1
X_11001_ net2399 net996 net337 VGND VGND VPWR VPWR _02745_ sky130_fd_sc_hd__mux2_1
XFILLER_120_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout850 net851 VGND VGND VPWR VPWR net850 sky130_fd_sc_hd__buf_12
Xfanout861 _05544_ VGND VGND VPWR VPWR net861 sky130_fd_sc_hd__clkbuf_1
Xfanout872 _05538_ VGND VGND VPWR VPWR net872 sky130_fd_sc_hd__clkbuf_2
Xfanout883 _05534_ VGND VGND VPWR VPWR net883 sky130_fd_sc_hd__clkbuf_2
Xfanout894 _05528_ VGND VGND VPWR VPWR net894 sky130_fd_sc_hd__clkbuf_2
XFILLER_18_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12952_ clknet_leaf_12_clk _01646_ VGND VGND VPWR VPWR data_array.data0\[13\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1070 data_array.data1\[6\]\[17\] VGND VGND VPWR VPWR net2721 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1081 tag_array.tag0\[0\]\[0\] VGND VGND VPWR VPWR net2732 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_133_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1092 data_array.data0\[3\]\[58\] VGND VGND VPWR VPWR net2743 sky130_fd_sc_hd__dlygate4sd3_1
X_11903_ clknet_leaf_244_clk _00711_ VGND VGND VPWR VPWR data_array.data0\[5\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
X_12883_ clknet_leaf_4_clk _01577_ VGND VGND VPWR VPWR data_array.data0\[12\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_61_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11834_ clknet_leaf_114_clk _00642_ VGND VGND VPWR VPWR data_array.data0\[7\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
X_11765_ clknet_leaf_38_clk _00573_ VGND VGND VPWR VPWR data_array.data0\[8\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_13504_ clknet_leaf_266_clk _02133_ VGND VGND VPWR VPWR data_array.data1\[0\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_10716_ net1110 net2855 net494 VGND VGND VPWR VPWR _02461_ sky130_fd_sc_hd__mux2_1
X_11696_ clknet_leaf_166_clk _00504_ VGND VGND VPWR VPWR tag_array.tag1\[15\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_14484_ clknet_leaf_165_clk _03107_ VGND VGND VPWR VPWR tag_array.dirty0\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_158_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13435_ clknet_leaf_20_clk _02065_ VGND VGND VPWR VPWR data_array.data1\[8\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
X_10647_ net1885 net874 net471 VGND VGND VPWR VPWR _02392_ sky130_fd_sc_hd__mux2_1
XFILLER_127_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload207 clknet_leaf_114_clk VGND VGND VPWR VPWR clkload207/X sky130_fd_sc_hd__clkbuf_4
XFILLER_9_189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload218 clknet_leaf_125_clk VGND VGND VPWR VPWR clkload218/Y sky130_fd_sc_hd__inv_6
Xrebuffer4 fsm.tag_out0\[0\] VGND VGND VPWR VPWR net1655 sky130_fd_sc_hd__dlygate4sd1_1
Xclkload229 clknet_leaf_157_clk VGND VGND VPWR VPWR clkload229/X sky130_fd_sc_hd__clkbuf_4
XFILLER_173_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13366_ clknet_leaf_165_clk _01996_ VGND VGND VPWR VPWR tag_array.tag0\[2\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_177_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10578_ net893 net2458 net454 VGND VGND VPWR VPWR _02323_ sky130_fd_sc_hd__mux2_1
XFILLER_127_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12317_ clknet_leaf_188_clk _01075_ VGND VGND VPWR VPWR tag_array.tag1\[12\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_177_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13297_ clknet_leaf_1_clk _01927_ VGND VGND VPWR VPWR data_array.data0\[10\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_114_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12248_ clknet_leaf_136_clk _01006_ VGND VGND VPWR VPWR tag_array.tag1\[14\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_131_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12179_ clknet_leaf_164_clk _00987_ VGND VGND VPWR VPWR tag_array.tag0\[14\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_95_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06740_ data_array.data0\[0\]\[0\] net1365 net1271 data_array.data0\[3\]\[0\] _04044_
+ VGND VGND VPWR VPWR _04045_ sky130_fd_sc_hd__a221o_1
XFILLER_95_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06671_ tag_array.tag1\[9\]\[19\] net1595 net1499 tag_array.tag1\[10\]\[19\] VGND
+ VGND VPWR VPWR _03982_ sky130_fd_sc_hd__a22o_1
X_08410_ net1124 _05509_ VGND VGND VPWR VPWR _05510_ sky130_fd_sc_hd__and2_1
X_05622_ fsm.tag_out1\[20\] VGND VGND VPWR VPWR _03144_ sky130_fd_sc_hd__inv_2
XFILLER_18_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09390_ net1104 net3461 net578 VGND VGND VPWR VPWR _01143_ sky130_fd_sc_hd__mux2_1
XFILLER_36_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_177_3761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08341_ net1124 _05463_ VGND VGND VPWR VPWR _05464_ sky130_fd_sc_hd__and2_1
XFILLER_178_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08272_ net807 _05416_ VGND VGND VPWR VPWR _05417_ sky130_fd_sc_hd__and2_4
XTAP_TAPCELL_ROW_15_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07223_ data_array.data0\[1\]\[44\] net1586 net1490 data_array.data0\[2\]\[44\] VGND
+ VGND VPWR VPWR _04484_ sky130_fd_sc_hd__a22o_1
XFILLER_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1080 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07154_ _04420_ _04421_ VGND VGND VPWR VPWR _00030_ sky130_fd_sc_hd__or2_1
X_06105_ data_array.rdata0\[20\] net1141 net1119 data_array.rdata1\[20\] VGND VGND
+ VPWR VPWR net275 sky130_fd_sc_hd__a22o_1
X_07085_ data_array.data0\[0\]\[31\] net1384 net1290 data_array.data0\[3\]\[31\] _04358_
+ VGND VGND VPWR VPWR _04359_ sky130_fd_sc_hd__a221o_1
X_06036_ fsm.tag_out0\[0\] net1121 _03481_ VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__a21o_1
XFILLER_133_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07987_ data_array.data1\[4\]\[49\] net1380 net1286 data_array.data1\[7\]\[49\] _05178_
+ VGND VGND VPWR VPWR _05179_ sky130_fd_sc_hd__a221o_1
XFILLER_41_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1043 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06938_ data_array.data0\[4\]\[18\] net1377 net1283 data_array.data0\[7\]\[18\] _04224_
+ VGND VGND VPWR VPWR _04225_ sky130_fd_sc_hd__a221o_1
X_09726_ net783 net3613 net676 VGND VGND VPWR VPWR _01478_ sky130_fd_sc_hd__mux2_1
XFILLER_41_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06869_ data_array.data0\[9\]\[12\] net1595 net1499 data_array.data0\[10\]\[12\]
+ VGND VGND VPWR VPWR _04162_ sky130_fd_sc_hd__a22o_1
X_09657_ net758 net3792 net614 VGND VGND VPWR VPWR _01409_ sky130_fd_sc_hd__mux2_1
XFILLER_83_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08608_ net791 net2808 net519 VGND VGND VPWR VPWR _00367_ sky130_fd_sc_hd__mux2_1
X_09588_ net998 net4063 net398 VGND VGND VPWR VPWR _01340_ sky130_fd_sc_hd__mux2_1
XFILLER_103_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08539_ net824 net815 net855 _05595_ VGND VGND VPWR VPWR _05597_ sky130_fd_sc_hd__or4_1
XFILLER_179_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11550_ clknet_leaf_140_clk _00358_ VGND VGND VPWR VPWR tag_array.tag1\[6\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_169_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10501_ net940 net3093 net350 VGND VGND VPWR VPWR _02246_ sky130_fd_sc_hd__mux2_1
XFILLER_184_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11481_ clknet_leaf_156_clk _00290_ VGND VGND VPWR VPWR tag_array.valid0\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_155_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13220_ clknet_leaf_252_clk _00116_ VGND VGND VPWR VPWR data_array.rdata1\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10432_ net2298 net924 net661 VGND VGND VPWR VPWR _02178_ sky130_fd_sc_hd__mux2_1
XFILLER_10_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13151_ clknet_leaf_134_clk _01845_ VGND VGND VPWR VPWR tag_array.tag1\[8\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_10363_ net749 net2564 net538 VGND VGND VPWR VPWR _02110_ sky130_fd_sc_hd__mux2_1
XFILLER_128_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12102_ clknet_leaf_75_clk _00910_ VGND VGND VPWR VPWR data_array.data1\[14\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
X_13082_ clknet_leaf_75_clk _01776_ VGND VGND VPWR VPWR data_array.data1\[13\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_112_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10294_ net2155 net985 net639 VGND VGND VPWR VPWR _02041_ sky130_fd_sc_hd__mux2_1
XFILLER_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12033_ clknet_leaf_49_clk _00841_ VGND VGND VPWR VPWR data_array.data0\[6\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout1601 net1603 VGND VGND VPWR VPWR net1601 sky130_fd_sc_hd__clkbuf_4
Xfanout1612 net1613 VGND VGND VPWR VPWR net1612 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_72_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1623 net1624 VGND VGND VPWR VPWR net1623 sky130_fd_sc_hd__buf_2
XFILLER_78_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1634 net1637 VGND VGND VPWR VPWR net1634 sky130_fd_sc_hd__buf_4
Xfanout1645 net98 VGND VGND VPWR VPWR net1645 sky130_fd_sc_hd__buf_4
XFILLER_66_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout680 net685 VGND VGND VPWR VPWR net680 sky130_fd_sc_hd__clkbuf_8
Xfanout691 net692 VGND VGND VPWR VPWR net691 sky130_fd_sc_hd__buf_4
X_13984_ clknet_leaf_91_clk _02613_ VGND VGND VPWR VPWR data_array.data1\[5\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_46_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12935_ clknet_leaf_234_clk _01629_ VGND VGND VPWR VPWR data_array.data0\[13\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12866_ clknet_leaf_10_clk _01560_ VGND VGND VPWR VPWR data_array.data0\[12\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_57_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11817_ clknet_leaf_59_clk _00625_ VGND VGND VPWR VPWR data_array.data0\[7\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_12797_ clknet_leaf_99_clk _01491_ VGND VGND VPWR VPWR tag_array.tag1\[10\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_155_3344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11748_ clknet_leaf_50_clk _00556_ VGND VGND VPWR VPWR data_array.data0\[8\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_147_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14467_ clknet_leaf_4_clk _03090_ VGND VGND VPWR VPWR data_array.data1\[7\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_146_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11679_ clknet_leaf_234_clk _00487_ VGND VGND VPWR VPWR tag_array.tag1\[1\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_13418_ clknet_leaf_77_clk _02048_ VGND VGND VPWR VPWR data_array.data1\[8\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_133_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14398_ clknet_leaf_76_clk _03021_ VGND VGND VPWR VPWR data_array.data1\[10\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_180_Right_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13349_ clknet_leaf_207_clk _01979_ VGND VGND VPWR VPWR data_array.data0\[10\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07910_ data_array.data1\[0\]\[42\] net1399 net1305 data_array.data1\[3\]\[42\] _05108_
+ VGND VGND VPWR VPWR _05109_ sky130_fd_sc_hd__a221o_1
Xhold2507 tag_array.tag1\[11\]\[23\] VGND VGND VPWR VPWR net4158 sky130_fd_sc_hd__dlygate4sd3_1
X_08890_ net945 net3162 net434 VGND VGND VPWR VPWR _00647_ sky130_fd_sc_hd__mux2_1
Xhold2518 data_array.data1\[10\]\[12\] VGND VGND VPWR VPWR net4169 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_25_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2529 data_array.data0\[7\]\[19\] VGND VGND VPWR VPWR net4180 sky130_fd_sc_hd__dlygate4sd3_1
X_07841_ data_array.data1\[13\]\[36\] net1606 net1510 data_array.data1\[14\]\[36\]
+ VGND VGND VPWR VPWR _05046_ sky130_fd_sc_hd__a22o_1
Xhold1806 lru_array.lru_mem\[8\] VGND VGND VPWR VPWR net3457 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1817 data_array.data0\[7\]\[8\] VGND VGND VPWR VPWR net3468 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1828 tag_array.tag0\[15\]\[0\] VGND VGND VPWR VPWR net3479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1839 data_array.data1\[5\]\[3\] VGND VGND VPWR VPWR net3490 sky130_fd_sc_hd__dlygate4sd3_1
X_07772_ data_array.data1\[8\]\[30\] net1393 net1299 data_array.data1\[11\]\[30\]
+ _04982_ VGND VGND VPWR VPWR _04983_ sky130_fd_sc_hd__a221o_1
XFILLER_84_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_179_3801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06723_ net1636 _04023_ _04027_ net1210 VGND VGND VPWR VPWR _04030_ sky130_fd_sc_hd__a22o_1
X_09511_ net785 net2833 net621 VGND VGND VPWR VPWR _01264_ sky130_fd_sc_hd__mux2_1
XFILLER_80_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09442_ net898 net3692 net578 VGND VGND VPWR VPWR _01195_ sky130_fd_sc_hd__mux2_1
X_06654_ tag_array.tag1\[8\]\[17\] net1421 net1327 tag_array.tag1\[11\]\[17\] _03966_
+ VGND VGND VPWR VPWR _03967_ sky130_fd_sc_hd__a221o_1
XFILLER_80_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09373_ net909 net3122 net403 VGND VGND VPWR VPWR _01126_ sky130_fd_sc_hd__mux2_1
XFILLER_12_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06585_ tag_array.tag1\[5\]\[11\] net1575 net1479 tag_array.tag1\[6\]\[11\] VGND
+ VGND VPWR VPWR _03904_ sky130_fd_sc_hd__a22o_1
XFILLER_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08324_ net2381 net1046 net689 VGND VGND VPWR VPWR _00237_ sky130_fd_sc_hd__mux2_1
XFILLER_71_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08255_ fsm.tag_out1\[20\] net816 net808 fsm.tag_out0\[20\] _05404_ VGND VGND VPWR
+ VPWR _05405_ sky130_fd_sc_hd__a221o_2
XFILLER_138_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07206_ data_array.data0\[0\]\[42\] net1388 net1294 data_array.data0\[3\]\[42\] _04468_
+ VGND VGND VPWR VPWR _04469_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_31_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08186_ net819 net2873 _05354_ VGND VGND VPWR VPWR _00195_ sky130_fd_sc_hd__mux2_1
XFILLER_174_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07137_ data_array.data0\[13\]\[36\] net1601 net1505 data_array.data0\[14\]\[36\]
+ VGND VGND VPWR VPWR _04406_ sky130_fd_sc_hd__a22o_1
XFILLER_119_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07068_ data_array.data0\[8\]\[30\] net1393 net1299 data_array.data0\[11\]\[30\]
+ _04342_ VGND VGND VPWR VPWR _04343_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_54_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput250 net250 VGND VGND VPWR VPWR mem_addr[28] sky130_fd_sc_hd__buf_2
Xoutput261 net261 VGND VGND VPWR VPWR mem_addr[9] sky130_fd_sc_hd__buf_2
X_06019_ net157 net1157 _03472_ _03473_ VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_54_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput272 net272 VGND VGND VPWR VPWR mem_wdata[18] sky130_fd_sc_hd__buf_2
Xoutput283 net283 VGND VGND VPWR VPWR mem_wdata[28] sky130_fd_sc_hd__buf_2
Xoutput294 net294 VGND VGND VPWR VPWR mem_wdata[38] sky130_fd_sc_hd__buf_2
XFILLER_181_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_50_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09709_ net752 net3761 net610 VGND VGND VPWR VPWR _01461_ sky130_fd_sc_hd__mux2_1
X_10981_ net1915 net1076 net337 VGND VGND VPWR VPWR _02725_ sky130_fd_sc_hd__mux2_1
XFILLER_16_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12720_ clknet_leaf_146_clk _01414_ VGND VGND VPWR VPWR tag_array.tag0\[7\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12651_ clknet_leaf_72_clk _01345_ VGND VGND VPWR VPWR data_array.data0\[15\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11602_ clknet_leaf_189_clk _00410_ VGND VGND VPWR VPWR tag_array.tag1\[4\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12582_ clknet_leaf_173_clk _01276_ VGND VGND VPWR VPWR tag_array.tag0\[10\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14321_ clknet_leaf_258_clk _02950_ VGND VGND VPWR VPWR data_array.data1\[11\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
X_11533_ clknet_leaf_152_clk _00341_ VGND VGND VPWR VPWR tag_array.valid0\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_183_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14252_ clknet_leaf_118_clk _02881_ VGND VGND VPWR VPWR data_array.data1\[12\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
X_11464_ clknet_leaf_3_clk _00274_ VGND VGND VPWR VPWR data_array.data0\[0\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_150_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13203_ clknet_leaf_122_clk _00098_ VGND VGND VPWR VPWR data_array.rdata1\[40\] sky130_fd_sc_hd__dfxtp_1
X_10415_ net1968 net994 net667 VGND VGND VPWR VPWR _02161_ sky130_fd_sc_hd__mux2_1
XFILLER_109_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14183_ clknet_leaf_37_clk _02812_ VGND VGND VPWR VPWR data_array.data0\[2\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_11395_ clknet_leaf_127_clk _00205_ VGND VGND VPWR VPWR tag_array.tag1\[7\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_111_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13134_ clknet_leaf_156_clk _01828_ VGND VGND VPWR VPWR tag_array.tag0\[3\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_10346_ net717 net4016 net592 VGND VGND VPWR VPWR _02093_ sky130_fd_sc_hd__mux2_1
XFILLER_180_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13065_ clknet_leaf_218_clk _01759_ VGND VGND VPWR VPWR data_array.data1\[13\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10277_ net1760 net1055 net639 VGND VGND VPWR VPWR _02024_ sky130_fd_sc_hd__mux2_1
Xfanout1420 net1421 VGND VGND VPWR VPWR net1420 sky130_fd_sc_hd__clkbuf_4
X_12016_ clknet_leaf_247_clk _00824_ VGND VGND VPWR VPWR data_array.data0\[6\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout1431 net1433 VGND VGND VPWR VPWR net1431 sky130_fd_sc_hd__clkbuf_4
XFILLER_94_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1442 net1443 VGND VGND VPWR VPWR net1442 sky130_fd_sc_hd__clkbuf_4
Xfanout1453 net1458 VGND VGND VPWR VPWR net1453 sky130_fd_sc_hd__buf_2
Xfanout1464 net1470 VGND VGND VPWR VPWR net1464 sky130_fd_sc_hd__buf_2
Xfanout1475 net1477 VGND VGND VPWR VPWR net1475 sky130_fd_sc_hd__clkbuf_2
Xfanout1486 net1495 VGND VGND VPWR VPWR net1486 sky130_fd_sc_hd__clkbuf_4
Xfanout1497 net1498 VGND VGND VPWR VPWR net1497 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13967_ clknet_leaf_82_clk _02596_ VGND VGND VPWR VPWR data_array.data1\[5\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_65_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12918_ clknet_leaf_22_clk _01612_ VGND VGND VPWR VPWR data_array.data0\[13\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_17_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13898_ clknet_leaf_215_clk _02527_ VGND VGND VPWR VPWR data_array.data1\[4\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12849_ clknet_leaf_249_clk _01543_ VGND VGND VPWR VPWR data_array.data0\[12\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_06370_ tag_array.tag0\[0\]\[16\] net1407 net1313 tag_array.tag0\[3\]\[16\] _03708_
+ VGND VGND VPWR VPWR _03709_ sky130_fd_sc_hd__a221o_1
XFILLER_159_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_170_3628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08040_ data_array.data1\[12\]\[54\] net1353 net1259 data_array.data1\[15\]\[54\]
+ _05226_ VGND VGND VPWR VPWR _05227_ sky130_fd_sc_hd__a221o_1
XFILLER_174_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold903 data_array.data0\[9\]\[24\] VGND VGND VPWR VPWR net2554 sky130_fd_sc_hd__dlygate4sd3_1
Xhold914 tag_array.tag1\[0\]\[7\] VGND VGND VPWR VPWR net2565 sky130_fd_sc_hd__dlygate4sd3_1
Xhold925 data_array.data1\[5\]\[36\] VGND VGND VPWR VPWR net2576 sky130_fd_sc_hd__dlygate4sd3_1
Xhold936 data_array.data1\[2\]\[59\] VGND VGND VPWR VPWR net2587 sky130_fd_sc_hd__dlygate4sd3_1
Xhold947 tag_array.tag1\[6\]\[4\] VGND VGND VPWR VPWR net2598 sky130_fd_sc_hd__dlygate4sd3_1
Xhold958 tag_array.tag0\[14\]\[21\] VGND VGND VPWR VPWR net2609 sky130_fd_sc_hd__dlygate4sd3_1
Xhold969 data_array.data1\[7\]\[40\] VGND VGND VPWR VPWR net2620 sky130_fd_sc_hd__dlygate4sd3_1
X_09991_ net866 net2923 net372 VGND VGND VPWR VPWR _01740_ sky130_fd_sc_hd__mux2_1
XFILLER_142_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08942_ net996 net3345 net427 VGND VGND VPWR VPWR _00698_ sky130_fd_sc_hd__mux2_1
Xhold2304 data_array.data0\[6\]\[21\] VGND VGND VPWR VPWR net3955 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2315 data_array.data0\[14\]\[17\] VGND VGND VPWR VPWR net3966 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2326 data_array.data0\[7\]\[3\] VGND VGND VPWR VPWR net3977 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2337 data_array.data0\[3\]\[27\] VGND VGND VPWR VPWR net3988 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2348 data_array.data1\[14\]\[39\] VGND VGND VPWR VPWR net3999 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1603 tag_array.tag1\[10\]\[0\] VGND VGND VPWR VPWR net3254 sky130_fd_sc_hd__dlygate4sd3_1
X_08873_ net1013 net2959 net440 VGND VGND VPWR VPWR _00630_ sky130_fd_sc_hd__mux2_1
Xhold1614 data_array.data1\[6\]\[62\] VGND VGND VPWR VPWR net3265 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2359 tag_array.tag1\[7\]\[17\] VGND VGND VPWR VPWR net4010 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1625 tag_array.tag0\[14\]\[0\] VGND VGND VPWR VPWR net3276 sky130_fd_sc_hd__dlygate4sd3_1
X_07824_ net1168 _05025_ _05029_ net1216 VGND VGND VPWR VPWR _05031_ sky130_fd_sc_hd__a22o_1
Xhold1636 tag_array.tag0\[1\]\[17\] VGND VGND VPWR VPWR net3287 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1647 data_array.data0\[3\]\[63\] VGND VGND VPWR VPWR net3298 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_659 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1658 tag_array.tag0\[0\]\[10\] VGND VGND VPWR VPWR net3309 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1669 data_array.data0\[13\]\[30\] VGND VGND VPWR VPWR net3320 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07755_ data_array.data1\[1\]\[28\] net1541 net1445 data_array.data1\[2\]\[28\] VGND
+ VGND VPWR VPWR _04968_ sky130_fd_sc_hd__a22o_1
X_06706_ tag_array.tag1\[1\]\[22\] net1552 net1456 tag_array.tag1\[2\]\[22\] VGND
+ VGND VPWR VPWR _04014_ sky130_fd_sc_hd__a22o_1
X_07686_ data_array.data1\[0\]\[22\] net1346 net1252 data_array.data1\[3\]\[22\] _04904_
+ VGND VGND VPWR VPWR _04905_ sky130_fd_sc_hd__a221o_1
X_09425_ net966 net2491 net586 VGND VGND VPWR VPWR _01178_ sky130_fd_sc_hd__mux2_1
X_06637_ _03950_ _03951_ VGND VGND VPWR VPWR _00162_ sky130_fd_sc_hd__or2_2
XFILLER_13_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06568_ tag_array.tag1\[0\]\[9\] net1418 net1324 tag_array.tag1\[3\]\[9\] _03888_
+ VGND VGND VPWR VPWR _03889_ sky130_fd_sc_hd__a221o_1
X_09356_ net977 net3091 net407 VGND VGND VPWR VPWR _01109_ sky130_fd_sc_hd__mux2_1
XFILLER_12_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08307_ net101 net36 net1640 VGND VGND VPWR VPWR _05441_ sky130_fd_sc_hd__mux2_1
X_09287_ net731 net4027 net561 VGND VGND VPWR VPWR _01041_ sky130_fd_sc_hd__mux2_1
X_06499_ tag_array.tag1\[13\]\[3\] net1561 net1465 tag_array.tag1\[14\]\[3\] VGND
+ VGND VPWR VPWR _03826_ sky130_fd_sc_hd__a22o_1
XFILLER_138_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_48 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08238_ net735 net3386 net799 VGND VGND VPWR VPWR _00210_ sky130_fd_sc_hd__mux2_1
XFILLER_181_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08169_ lru_array.lru_mem\[5\] net1563 net1467 lru_array.lru_mem\[6\] VGND VGND VPWR
+ VPWR _05344_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_91_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10200_ net1006 net3721 net355 VGND VGND VPWR VPWR _01947_ sky130_fd_sc_hd__mux2_1
XFILLER_118_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11180_ net1055 net3110 net655 VGND VGND VPWR VPWR _02923_ sky130_fd_sc_hd__mux2_1
XFILLER_69_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10131_ net1022 net3826 net363 VGND VGND VPWR VPWR _01879_ sky130_fd_sc_hd__mux2_1
XFILLER_133_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10062_ net776 net3835 net599 VGND VGND VPWR VPWR _01811_ sky130_fd_sc_hd__mux2_1
XFILLER_0_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2860 data_array.data1\[9\]\[28\] VGND VGND VPWR VPWR net4511 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2871 data_array.data1\[12\]\[9\] VGND VGND VPWR VPWR net4522 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2882 data_array.data0\[5\]\[31\] VGND VGND VPWR VPWR net4533 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2893 tag_array.tag0\[0\]\[20\] VGND VGND VPWR VPWR net4544 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13821_ clknet_leaf_8_clk _02450_ VGND VGND VPWR VPWR data_array.data1\[2\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13752_ clknet_leaf_75_clk _02381_ VGND VGND VPWR VPWR data_array.data1\[1\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_141_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10964_ net886 net2845 net527 VGND VGND VPWR VPWR _02709_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_67_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12703_ clknet_leaf_156_clk _01397_ VGND VGND VPWR VPWR tag_array.tag0\[8\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_44_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_104_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13683_ clknet_leaf_43_clk _02312_ VGND VGND VPWR VPWR data_array.data1\[15\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
X_10895_ net906 net4241 net514 VGND VGND VPWR VPWR _02640_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_84_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12634_ clknet_leaf_222_clk _01328_ VGND VGND VPWR VPWR data_array.data0\[15\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_169_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12565_ clknet_leaf_185_clk _01259_ VGND VGND VPWR VPWR tag_array.tag0\[11\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14304_ clknet_leaf_89_clk _02933_ VGND VGND VPWR VPWR data_array.data1\[11\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11516_ clknet_leaf_99_clk _00324_ VGND VGND VPWR VPWR tag_array.tag1\[9\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_12496_ clknet_leaf_76_clk _01190_ VGND VGND VPWR VPWR data_array.data1\[9\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_157_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_44_Left_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14235_ clknet_leaf_67_clk _02864_ VGND VGND VPWR VPWR data_array.data1\[12\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_171_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11447_ clknet_leaf_113_clk _00257_ VGND VGND VPWR VPWR data_array.data0\[0\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_125_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11378_ net819 net3246 _05581_ VGND VGND VPWR VPWR _03121_ sky130_fd_sc_hd__mux2_1
XFILLER_98_504 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14166_ clknet_leaf_49_clk _02795_ VGND VGND VPWR VPWR data_array.data0\[2\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_125_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13117_ clknet_leaf_177_clk _01811_ VGND VGND VPWR VPWR tag_array.tag0\[3\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_10329_ net784 net4550 net591 VGND VGND VPWR VPWR _02076_ sky130_fd_sc_hd__mux2_1
XFILLER_98_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14097_ clknet_leaf_62_clk _02726_ VGND VGND VPWR VPWR data_array.data0\[1\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_13048_ clknet_leaf_224_clk _01742_ VGND VGND VPWR VPWR data_array.data0\[3\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_38_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1250 net1251 VGND VGND VPWR VPWR net1250 sky130_fd_sc_hd__clkbuf_4
Xfanout1261 net1270 VGND VGND VPWR VPWR net1261 sky130_fd_sc_hd__buf_2
X_05870_ data_array.rdata0\[13\] net848 net1145 VGND VGND VPWR VPWR _03374_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_163_3487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1272 net1273 VGND VGND VPWR VPWR net1272 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_163_3498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1283 net1284 VGND VGND VPWR VPWR net1283 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_1_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1294 net1306 VGND VGND VPWR VPWR net1294 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_1_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_53_Left_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07540_ data_array.data1\[9\]\[9\] net1581 net1485 data_array.data1\[10\]\[9\] VGND
+ VGND VPWR VPWR _04772_ sky130_fd_sc_hd__a22o_1
XFILLER_179_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07471_ net1190 _04703_ _04707_ net1616 VGND VGND VPWR VPWR _04710_ sky130_fd_sc_hd__a22o_1
XFILLER_90_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06422_ tag_array.tag0\[9\]\[21\] net1600 net1504 tag_array.tag0\[10\]\[21\] VGND
+ VGND VPWR VPWR _03756_ sky130_fd_sc_hd__a22o_1
X_09210_ net738 net2525 net631 VGND VGND VPWR VPWR _00964_ sky130_fd_sc_hd__mux2_1
XFILLER_148_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09141_ net978 net4475 net574 VGND VGND VPWR VPWR _00895_ sky130_fd_sc_hd__mux2_1
X_06353_ tag_array.tag0\[12\]\[15\] net1402 net1308 tag_array.tag0\[15\]\[15\] _03692_
+ VGND VGND VPWR VPWR _03693_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_62_Left_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09072_ net996 net2480 net411 VGND VGND VPWR VPWR _00826_ sky130_fd_sc_hd__mux2_1
X_06284_ net1230 _03625_ _03629_ net1182 VGND VGND VPWR VPWR _03631_ sky130_fd_sc_hd__a22o_1
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08023_ _05210_ _05211_ VGND VGND VPWR VPWR _00111_ sky130_fd_sc_hd__or2_1
Xhold700 tag_array.tag1\[9\]\[2\] VGND VGND VPWR VPWR net2351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold711 data_array.data1\[15\]\[23\] VGND VGND VPWR VPWR net2362 sky130_fd_sc_hd__dlygate4sd3_1
Xhold722 data_array.data1\[8\]\[36\] VGND VGND VPWR VPWR net2373 sky130_fd_sc_hd__dlygate4sd3_1
Xhold733 data_array.data0\[0\]\[13\] VGND VGND VPWR VPWR net2384 sky130_fd_sc_hd__dlygate4sd3_1
Xhold744 tag_array.tag1\[15\]\[2\] VGND VGND VPWR VPWR net2395 sky130_fd_sc_hd__dlygate4sd3_1
Xhold755 data_array.data1\[1\]\[40\] VGND VGND VPWR VPWR net2406 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold766 tag_array.tag0\[14\]\[2\] VGND VGND VPWR VPWR net2417 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold777 data_array.data1\[4\]\[31\] VGND VGND VPWR VPWR net2428 sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 data_array.data1\[3\]\[60\] VGND VGND VPWR VPWR net2439 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09974_ net932 net3250 _03127_ VGND VGND VPWR VPWR _01723_ sky130_fd_sc_hd__mux2_1
Xhold799 data_array.data0\[13\]\[21\] VGND VGND VPWR VPWR net2450 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2101 tag_array.tag0\[5\]\[16\] VGND VGND VPWR VPWR net3752 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2112 data_array.data1\[11\]\[12\] VGND VGND VPWR VPWR net3763 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2123 data_array.data1\[11\]\[35\] VGND VGND VPWR VPWR net3774 sky130_fd_sc_hd__dlygate4sd3_1
X_08925_ net1064 net2531 net431 VGND VGND VPWR VPWR _00681_ sky130_fd_sc_hd__mux2_1
Xhold2134 tag_array.tag0\[12\]\[10\] VGND VGND VPWR VPWR net3785 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2145 tag_array.tag1\[11\]\[24\] VGND VGND VPWR VPWR net3796 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1400 data_array.data0\[2\]\[43\] VGND VGND VPWR VPWR net3051 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1411 data_array.data0\[14\]\[41\] VGND VGND VPWR VPWR net3062 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_71_Left_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2156 tag_array.tag0\[4\]\[8\] VGND VGND VPWR VPWR net3807 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1422 data_array.data1\[12\]\[42\] VGND VGND VPWR VPWR net3073 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2167 data_array.data0\[10\]\[23\] VGND VGND VPWR VPWR net3818 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1433 tag_array.dirty1\[13\] VGND VGND VPWR VPWR net3084 sky130_fd_sc_hd__dlygate4sd3_1
X_08856_ net1080 net2338 net440 VGND VGND VPWR VPWR _00613_ sky130_fd_sc_hd__mux2_1
Xhold2178 data_array.data0\[10\]\[28\] VGND VGND VPWR VPWR net3829 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2189 tag_array.tag0\[3\]\[14\] VGND VGND VPWR VPWR net3840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1444 tag_array.tag0\[9\]\[24\] VGND VGND VPWR VPWR net3095 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1455 tag_array.tag0\[4\]\[22\] VGND VGND VPWR VPWR net3106 sky130_fd_sc_hd__dlygate4sd3_1
X_07807_ data_array.data1\[0\]\[33\] net1397 net1303 data_array.data1\[3\]\[33\] _05014_
+ VGND VGND VPWR VPWR _05015_ sky130_fd_sc_hd__a221o_1
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1466 tag_array.tag0\[8\]\[3\] VGND VGND VPWR VPWR net3117 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1477 data_array.data0\[5\]\[18\] VGND VGND VPWR VPWR net3128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1488 data_array.data1\[3\]\[38\] VGND VGND VPWR VPWR net3139 sky130_fd_sc_hd__dlygate4sd3_1
X_05999_ data_array.rdata0\[56\] net853 net1146 VGND VGND VPWR VPWR _03460_ sky130_fd_sc_hd__o21a_1
X_08787_ net2222 net1097 net446 VGND VGND VPWR VPWR _00545_ sky130_fd_sc_hd__mux2_1
Xhold1499 data_array.data0\[14\]\[32\] VGND VGND VPWR VPWR net3150 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_49_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07738_ data_array.data1\[9\]\[27\] net1547 net1451 data_array.data1\[10\]\[27\]
+ VGND VGND VPWR VPWR _04952_ sky130_fd_sc_hd__a22o_1
XFILLER_164_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07669_ net1210 _04883_ _04887_ net1636 VGND VGND VPWR VPWR _04890_ sky130_fd_sc_hd__a22o_1
XFILLER_13_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09408_ net1035 net3380 net586 VGND VGND VPWR VPWR _01161_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10680_ net3184 net997 net479 VGND VGND VPWR VPWR _02425_ sky130_fd_sc_hd__mux2_1
XFILLER_179_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_80_Left_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09339_ net1046 net3493 net404 VGND VGND VPWR VPWR _01092_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_109_Right_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12350_ clknet_leaf_257_clk _00025_ VGND VGND VPWR VPWR data_array.rdata0\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_181_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11301_ net1090 net3065 net799 VGND VGND VPWR VPWR _03044_ sky130_fd_sc_hd__mux2_1
X_12281_ clknet_leaf_134_clk _01039_ VGND VGND VPWR VPWR tag_array.tag1\[13\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_14020_ clknet_leaf_120_clk _02649_ VGND VGND VPWR VPWR data_array.data1\[5\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
X_11232_ net1101 net4332 net674 VGND VGND VPWR VPWR _02975_ sky130_fd_sc_hd__mux2_1
XFILLER_5_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11163_ net865 net3048 net545 VGND VGND VPWR VPWR _02906_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10114_ net1089 net4128 net364 VGND VGND VPWR VPWR _01862_ sky130_fd_sc_hd__mux2_1
XFILLER_171_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11094_ net2685 net884 net329 VGND VGND VPWR VPWR _02837_ sky130_fd_sc_hd__mux2_1
XFILLER_110_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_145_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10045_ net906 net2772 net554 VGND VGND VPWR VPWR _01794_ sky130_fd_sc_hd__mux2_1
XFILLER_102_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold60 tag_array.valid0\[11\] VGND VGND VPWR VPWR net1711 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_69_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold71 tag_array.valid0\[0\] VGND VGND VPWR VPWR net1722 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 tag_array.tag1\[2\]\[16\] VGND VGND VPWR VPWR net1733 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2690 data_array.data0\[6\]\[43\] VGND VGND VPWR VPWR net4341 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold93 data_array.data1\[4\]\[43\] VGND VGND VPWR VPWR net1744 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_21_1041 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13804_ clknet_leaf_85_clk _02433_ VGND VGND VPWR VPWR data_array.data1\[2\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_91_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11996_ clknet_leaf_270_clk _00804_ VGND VGND VPWR VPWR data_array.data0\[6\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13735_ clknet_leaf_41_clk _02364_ VGND VGND VPWR VPWR data_array.data1\[1\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_10947_ net953 net4096 net527 VGND VGND VPWR VPWR _02692_ sky130_fd_sc_hd__mux2_1
XFILLER_45_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13666_ clknet_leaf_255_clk _02295_ VGND VGND VPWR VPWR data_array.data1\[15\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_10878_ net974 net2982 net515 VGND VGND VPWR VPWR _02623_ sky130_fd_sc_hd__mux2_1
X_12617_ clknet_leaf_186_clk _01311_ VGND VGND VPWR VPWR tag_array.tag0\[0\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_84_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13597_ clknet_leaf_22_clk _02226_ VGND VGND VPWR VPWR data_array.data0\[9\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_4_14_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_14_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_157_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12548_ clknet_leaf_147_clk _01242_ VGND VGND VPWR VPWR tag_array.tag0\[11\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_145_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_2 _00024_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12479_ clknet_leaf_37_clk _01173_ VGND VGND VPWR VPWR data_array.data1\[9\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14218_ clknet_leaf_251_clk _02847_ VGND VGND VPWR VPWR data_array.data1\[12\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_802 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_165_3527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14149_ clknet_leaf_206_clk _02778_ VGND VGND VPWR VPWR data_array.data0\[1\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout509 net512 VGND VGND VPWR VPWR net509 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_165_3538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_182_3852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06971_ data_array.data0\[0\]\[21\] net1366 net1272 data_array.data0\[3\]\[21\] _04254_
+ VGND VGND VPWR VPWR _04255_ sky130_fd_sc_hd__a221o_1
XFILLER_100_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_182_3863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08710_ net2055 net782 net474 VGND VGND VPWR VPWR _00469_ sky130_fd_sc_hd__mux2_1
XFILLER_140_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05922_ data_array.rdata1\[30\] net832 net841 VGND VGND VPWR VPWR _03409_ sky130_fd_sc_hd__a21o_1
X_09690_ net726 net3752 net606 VGND VGND VPWR VPWR _01442_ sky130_fd_sc_hd__mux2_1
XFILLER_67_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1080 net1081 VGND VGND VPWR VPWR net1080 sky130_fd_sc_hd__clkbuf_2
X_05853_ data_array.rdata1\[7\] net834 net843 VGND VGND VPWR VPWR _03363_ sky130_fd_sc_hd__a21o_1
Xfanout1091 _05430_ VGND VGND VPWR VPWR net1091 sky130_fd_sc_hd__dlymetal6s2s_1
X_08641_ net3001 net759 net511 VGND VGND VPWR VPWR _00400_ sky130_fd_sc_hd__mux2_1
XFILLER_82_724 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08572_ net812 _05583_ VGND VGND VPWR VPWR _05601_ sky130_fd_sc_hd__nand2_2
X_05784_ net2 fsm.tag_out1\[3\] VGND VGND VPWR VPWR _03301_ sky130_fd_sc_hd__and2b_1
X_07523_ data_array.data1\[12\]\[7\] net1398 net1304 data_array.data1\[15\]\[7\] _04756_
+ VGND VGND VPWR VPWR _04757_ sky130_fd_sc_hd__a221o_1
XFILLER_35_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07454_ data_array.data1\[1\]\[1\] net1520 net1424 data_array.data1\[2\]\[1\] VGND
+ VGND VPWR VPWR _04694_ sky130_fd_sc_hd__a22o_1
X_06405_ net1230 _03735_ _03739_ net1181 VGND VGND VPWR VPWR _03741_ sky130_fd_sc_hd__a22o_1
X_07385_ _04630_ _04631_ VGND VGND VPWR VPWR _00053_ sky130_fd_sc_hd__or2_1
XFILLER_109_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09124_ net1045 net3107 net570 VGND VGND VPWR VPWR _00878_ sky130_fd_sc_hd__mux2_1
XFILLER_109_918 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06336_ tag_array.tag0\[5\]\[13\] net1608 net1512 tag_array.tag0\[6\]\[13\] VGND
+ VGND VPWR VPWR _03678_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_40_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09055_ net1065 net4297 net415 VGND VGND VPWR VPWR _00809_ sky130_fd_sc_hd__mux2_1
X_06267_ tag_array.tag0\[0\]\[7\] net1418 net1324 tag_array.tag0\[3\]\[7\] _03614_
+ VGND VGND VPWR VPWR _03615_ sky130_fd_sc_hd__a221o_1
X_08006_ data_array.data1\[9\]\[51\] net1522 net1426 data_array.data1\[10\]\[51\]
+ VGND VGND VPWR VPWR _05196_ sky130_fd_sc_hd__a22o_1
Xhold530 data_array.data1\[4\]\[33\] VGND VGND VPWR VPWR net2181 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_163_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06198_ tag_array.tag0\[9\]\[1\] net1593 net1497 tag_array.tag0\[10\]\[1\] VGND VGND
+ VPWR VPWR _03552_ sky130_fd_sc_hd__a22o_1
Xhold541 data_array.data1\[0\]\[11\] VGND VGND VPWR VPWR net2192 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold552 data_array.data1\[1\]\[23\] VGND VGND VPWR VPWR net2203 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold563 tag_array.tag1\[8\]\[17\] VGND VGND VPWR VPWR net2214 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_173_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold574 data_array.data1\[1\]\[27\] VGND VGND VPWR VPWR net2225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold585 data_array.data1\[7\]\[63\] VGND VGND VPWR VPWR net2236 sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 data_array.data1\[1\]\[62\] VGND VGND VPWR VPWR net2247 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09957_ net1002 net3988 net373 VGND VGND VPWR VPWR _01706_ sky130_fd_sc_hd__mux2_1
X_08908_ net872 net4085 net438 VGND VGND VPWR VPWR _00665_ sky130_fd_sc_hd__mux2_1
X_09888_ net916 net2602 net383 VGND VGND VPWR VPWR _01638_ sky130_fd_sc_hd__mux2_1
Xhold1230 data_array.data0\[9\]\[46\] VGND VGND VPWR VPWR net2881 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1241 data_array.data1\[12\]\[30\] VGND VGND VPWR VPWR net2892 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_86_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1252 data_array.data0\[5\]\[46\] VGND VGND VPWR VPWR net2903 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_86_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08839_ net1943 net888 net443 VGND VGND VPWR VPWR _00597_ sky130_fd_sc_hd__mux2_1
Xhold1263 tag_array.tag0\[0\]\[14\] VGND VGND VPWR VPWR net2914 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1274 data_array.data0\[9\]\[25\] VGND VGND VPWR VPWR net2925 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1285 data_array.data1\[3\]\[22\] VGND VGND VPWR VPWR net2936 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1296 data_array.data1\[0\]\[33\] VGND VGND VPWR VPWR net2947 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_223 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11850_ clknet_leaf_208_clk _00658_ VGND VGND VPWR VPWR data_array.data0\[7\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_167_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10801_ net2741 net1024 net506 VGND VGND VPWR VPWR _02546_ sky130_fd_sc_hd__mux2_1
XFILLER_14_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ clknet_leaf_92_clk _00589_ VGND VGND VPWR VPWR data_array.data0\[8\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
X_13520_ clknet_leaf_253_clk _02149_ VGND VGND VPWR VPWR data_array.data1\[0\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_10732_ net1044 net4103 net493 VGND VGND VPWR VPWR _02477_ sky130_fd_sc_hd__mux2_1
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13451_ clknet_leaf_142_clk _02081_ VGND VGND VPWR VPWR tag_array.tag0\[1\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_10663_ net1811 net1067 net483 VGND VGND VPWR VPWR _02408_ sky130_fd_sc_hd__mux2_1
X_12402_ clknet_leaf_127_clk _01096_ VGND VGND VPWR VPWR data_array.data0\[14\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_13382_ clknet_leaf_251_clk _02012_ VGND VGND VPWR VPWR data_array.data1\[8\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_10594_ net1959 net1086 net466 VGND VGND VPWR VPWR _02339_ sky130_fd_sc_hd__mux2_1
XFILLER_51_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12333_ clknet_leaf_65_clk _00006_ VGND VGND VPWR VPWR data_array.rdata0\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12264_ clknet_leaf_103_clk _01022_ VGND VGND VPWR VPWR tag_array.tag1\[14\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_118_Left_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14003_ clknet_leaf_44_clk _02632_ VGND VGND VPWR VPWR data_array.data1\[5\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
X_11215_ net914 net3671 net655 VGND VGND VPWR VPWR _02958_ sky130_fd_sc_hd__mux2_1
XFILLER_141_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12195_ clknet_leaf_183_clk _00148_ VGND VGND VPWR VPWR fsm.tag_out0\[2\] sky130_fd_sc_hd__dfxtp_2
X_11146_ net935 net2585 net550 VGND VGND VPWR VPWR _02889_ sky130_fd_sc_hd__mux2_1
XFILLER_96_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11077_ net2515 net954 net332 VGND VGND VPWR VPWR _02820_ sky130_fd_sc_hd__mux2_1
XFILLER_163_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput150 mem_rdata[56] VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_160_3435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput161 mem_rdata[8] VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_160_3446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10028_ net975 net2499 net556 VGND VGND VPWR VPWR _01777_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_196_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_196_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_36_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_127_Left_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11979_ clknet_leaf_3_clk _00787_ VGND VGND VPWR VPWR data_array.data0\[4\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
X_13718_ clknet_leaf_47_clk _02347_ VGND VGND VPWR VPWR data_array.data1\[1\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_952 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_3397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13649_ clknet_leaf_57_clk _02278_ VGND VGND VPWR VPWR data_array.data1\[15\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_164_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07170_ data_array.data0\[13\]\[39\] net1541 net1445 data_array.data0\[14\]\[39\]
+ VGND VGND VPWR VPWR _04436_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_119_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06121_ data_array.rdata0\[36\] net1141 net1119 data_array.rdata1\[36\] VGND VGND
+ VPWR VPWR net292 sky130_fd_sc_hd__a22o_1
XFILLER_117_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_120_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_120_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_136_Left_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06052_ fsm.tag_out0\[8\] net1122 _03489_ VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_10_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_184_3903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_184_3914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_1074 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09811_ net965 net2601 net392 VGND VGND VPWR VPWR _01562_ sky130_fd_sc_hd__mux2_1
Xfanout328 net332 VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__buf_4
XFILLER_154_1066 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout339 net340 VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__clkbuf_4
XFILLER_101_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09742_ net719 net2285 net679 VGND VGND VPWR VPWR _01494_ sky130_fd_sc_hd__mux2_1
X_06954_ net1204 _04233_ _04237_ net1630 VGND VGND VPWR VPWR _04240_ sky130_fd_sc_hd__a22o_1
X_05905_ net115 net1155 _03396_ _03397_ VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__a22o_1
X_09673_ net696 net4527 net614 VGND VGND VPWR VPWR _01425_ sky130_fd_sc_hd__mux2_1
X_06885_ data_array.data0\[8\]\[13\] net1361 net1267 data_array.data0\[11\]\[13\]
+ _04176_ VGND VGND VPWR VPWR _04177_ sky130_fd_sc_hd__a221o_1
XFILLER_55_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_187_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_187_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_145_Left_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08624_ net729 net2724 net523 VGND VGND VPWR VPWR _00383_ sky130_fd_sc_hd__mux2_1
X_05836_ net110 net1150 _03350_ _03351_ VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__a22o_1
XFILLER_70_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08555_ net734 net3936 net584 VGND VGND VPWR VPWR _00323_ sky130_fd_sc_hd__mux2_1
X_05767_ _03276_ _03281_ _03282_ _03283_ VGND VGND VPWR VPWR _03284_ sky130_fd_sc_hd__or4_1
XFILLER_23_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07506_ _04740_ _04741_ VGND VGND VPWR VPWR _00119_ sky130_fd_sc_hd__or2_1
XFILLER_52_16 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08486_ net1273 net1173 net811 net1708 VGND VGND VPWR VPWR _00291_ sky130_fd_sc_hd__a31o_1
X_05698_ net18 _03145_ _03155_ _03209_ VGND VGND VPWR VPWR _03215_ sky130_fd_sc_hd__a211o_1
XFILLER_168_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07437_ data_array.data0\[0\]\[63\] net1358 net1264 data_array.data0\[3\]\[63\] _04678_
+ VGND VGND VPWR VPWR _04679_ sky130_fd_sc_hd__a221o_1
XFILLER_10_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07368_ data_array.data0\[9\]\[57\] net1555 net1459 data_array.data0\[10\]\[57\]
+ VGND VGND VPWR VPWR _04616_ sky130_fd_sc_hd__a22o_1
X_09107_ net856 net3180 net413 VGND VGND VPWR VPWR _00861_ sky130_fd_sc_hd__mux2_1
XFILLER_182_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06319_ tag_array.tag0\[9\]\[12\] net1597 net1501 tag_array.tag0\[10\]\[12\] VGND
+ VGND VPWR VPWR _03662_ sky130_fd_sc_hd__a22o_1
X_07299_ data_array.data0\[12\]\[51\] net1332 net1238 data_array.data0\[15\]\[51\]
+ _04552_ VGND VGND VPWR VPWR _04553_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_111_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_111_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_184_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09038_ net2167 net872 net422 VGND VGND VPWR VPWR _00793_ sky130_fd_sc_hd__mux2_1
XFILLER_163_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold360 data_array.data1\[8\]\[21\] VGND VGND VPWR VPWR net2011 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold371 data_array.data1\[4\]\[39\] VGND VGND VPWR VPWR net2022 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold382 data_array.data1\[4\]\[18\] VGND VGND VPWR VPWR net2033 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold393 data_array.data1\[0\]\[48\] VGND VGND VPWR VPWR net2044 sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ net2730 net1002 net339 VGND VGND VPWR VPWR _02744_ sky130_fd_sc_hd__mux2_1
XFILLER_105_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout840 net844 VGND VGND VPWR VPWR net840 sky130_fd_sc_hd__buf_6
Xfanout851 net852 VGND VGND VPWR VPWR net851 sky130_fd_sc_hd__buf_12
Xfanout862 _05544_ VGND VGND VPWR VPWR net862 sky130_fd_sc_hd__clkbuf_2
Xfanout873 _05538_ VGND VGND VPWR VPWR net873 sky130_fd_sc_hd__clkbuf_1
Xfanout884 _05532_ VGND VGND VPWR VPWR net884 sky130_fd_sc_hd__clkbuf_2
XFILLER_19_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout895 _05528_ VGND VGND VPWR VPWR net895 sky130_fd_sc_hd__buf_1
X_12951_ clknet_leaf_16_clk _01645_ VGND VGND VPWR VPWR data_array.data0\[13\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_178_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_178_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_19_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1060 data_array.data0\[0\]\[7\] VGND VGND VPWR VPWR net2711 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1071 data_array.data1\[13\]\[50\] VGND VGND VPWR VPWR net2722 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11902_ clknet_leaf_109_clk _00710_ VGND VGND VPWR VPWR data_array.data0\[5\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_46_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1082 tag_array.tag0\[11\]\[12\] VGND VGND VPWR VPWR net2733 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12882_ clknet_leaf_25_clk _01576_ VGND VGND VPWR VPWR data_array.data0\[12\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1093 tag_array.tag1\[2\]\[11\] VGND VGND VPWR VPWR net2744 sky130_fd_sc_hd__dlygate4sd3_1
X_11833_ clknet_leaf_242_clk _00641_ VGND VGND VPWR VPWR data_array.data0\[7\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11764_ clknet_leaf_69_clk _00572_ VGND VGND VPWR VPWR data_array.data0\[8\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_159_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_161_Right_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13503_ clknet_leaf_174_clk _02132_ VGND VGND VPWR VPWR data_array.data1\[0\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_10715_ net1788 net858 net481 VGND VGND VPWR VPWR _02460_ sky130_fd_sc_hd__mux2_1
X_14483_ clknet_leaf_101_clk _03106_ VGND VGND VPWR VPWR tag_array.dirty0\[2\] sky130_fd_sc_hd__dfxtp_1
X_11695_ clknet_leaf_33_clk _00503_ VGND VGND VPWR VPWR tag_array.tag1\[15\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_13434_ clknet_leaf_215_clk _02064_ VGND VGND VPWR VPWR data_array.data1\[8\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
X_10646_ net2077 net878 net470 VGND VGND VPWR VPWR _02391_ sky130_fd_sc_hd__mux2_1
Xclkload208 clknet_leaf_115_clk VGND VGND VPWR VPWR clkload208/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_158_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload219 clknet_leaf_126_clk VGND VGND VPWR VPWR clkload219/Y sky130_fd_sc_hd__clkinv_8
Xrebuffer5 fsm.tag_out0\[0\] VGND VGND VPWR VPWR net1656 sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_102_clk clknet_5_24__leaf_clk VGND VGND VPWR VPWR clknet_leaf_102_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13365_ clknet_leaf_105_clk _01995_ VGND VGND VPWR VPWR tag_array.tag0\[2\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_158_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10577_ net898 net4493 net453 VGND VGND VPWR VPWR _02322_ sky130_fd_sc_hd__mux2_1
XFILLER_177_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12316_ clknet_leaf_130_clk _01074_ VGND VGND VPWR VPWR tag_array.tag1\[12\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_155_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13296_ clknet_leaf_205_clk _01926_ VGND VGND VPWR VPWR data_array.data0\[10\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12247_ clknet_leaf_194_clk _01005_ VGND VGND VPWR VPWR tag_array.tag1\[14\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_131_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12178_ clknet_leaf_107_clk _00986_ VGND VGND VPWR VPWR tag_array.tag0\[14\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_11129_ net1001 net3088 net542 VGND VGND VPWR VPWR _02872_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_169_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_169_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_114_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06670_ _03980_ _03981_ VGND VGND VPWR VPWR _00165_ sky130_fd_sc_hd__or2_1
XFILLER_64_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05621_ net20 VGND VGND VPWR VPWR _03143_ sky130_fd_sc_hd__inv_2
XFILLER_184_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_177_3762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08340_ net113 net48 net1638 VGND VGND VPWR VPWR _05463_ sky130_fd_sc_hd__mux2_1
XFILLER_32_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08271_ _03514_ _03519_ VGND VGND VPWR VPWR _05416_ sky130_fd_sc_hd__nor2_1
XFILLER_178_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07222_ data_array.data0\[8\]\[44\] net1399 net1305 data_array.data0\[11\]\[44\]
+ _04482_ VGND VGND VPWR VPWR _04483_ sky130_fd_sc_hd__a221o_1
XFILLER_121_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07153_ net1218 _04415_ _04419_ net1170 VGND VGND VPWR VPWR _04421_ sky130_fd_sc_hd__a22o_1
XFILLER_121_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06104_ data_array.rdata0\[19\] net1139 net1115 data_array.rdata1\[19\] VGND VGND
+ VPWR VPWR net273 sky130_fd_sc_hd__a22o_1
XFILLER_118_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07084_ data_array.data0\[1\]\[31\] net1576 net1480 data_array.data0\[2\]\[31\] VGND
+ VGND VPWR VPWR _04358_ sky130_fd_sc_hd__a22o_1
XFILLER_118_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06035_ net1161 net30 fsm.tag_out1\[0\] net1132 VGND VGND VPWR VPWR _03481_ sky130_fd_sc_hd__a22o_1
XFILLER_114_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_5_28__f_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_5_28__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_35_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07986_ data_array.data1\[5\]\[49\] net1571 net1475 data_array.data1\[6\]\[49\] VGND
+ VGND VPWR VPWR _05178_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09725_ net786 net4616 net675 VGND VGND VPWR VPWR _01477_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06937_ data_array.data0\[5\]\[18\] net1567 net1471 data_array.data0\[6\]\[18\] VGND
+ VGND VPWR VPWR _04224_ sky130_fd_sc_hd__a22o_1
XFILLER_41_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09656_ net762 net4610 net614 VGND VGND VPWR VPWR _01408_ sky130_fd_sc_hd__mux2_1
X_06868_ _04160_ _04161_ VGND VGND VPWR VPWR _00002_ sky130_fd_sc_hd__or2_1
X_08607_ net694 net3768 net529 VGND VGND VPWR VPWR _00366_ sky130_fd_sc_hd__mux2_1
XFILLER_82_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_05819_ _03251_ _03263_ _03266_ _03270_ VGND VGND VPWR VPWR _03336_ sky130_fd_sc_hd__or4_1
X_09587_ net1002 net3210 net397 VGND VGND VPWR VPWR _01339_ sky130_fd_sc_hd__mux2_1
X_06799_ data_array.data0\[4\]\[5\] net1354 net1260 data_array.data0\[7\]\[5\] _04098_
+ VGND VGND VPWR VPWR _04099_ sky130_fd_sc_hd__a221o_1
XFILLER_179_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08538_ net825 _05595_ VGND VGND VPWR VPWR _05596_ sky130_fd_sc_hd__or2_1
XFILLER_11_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08469_ net812 _05416_ VGND VGND VPWR VPWR _05549_ sky130_fd_sc_hd__and2_2
X_10500_ net946 net3219 net345 VGND VGND VPWR VPWR _02245_ sky130_fd_sc_hd__mux2_1
XFILLER_128_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11480_ clknet_leaf_173_clk _00289_ VGND VGND VPWR VPWR tag_array.valid1\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_98_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10431_ net2009 net930 net663 VGND VGND VPWR VPWR _02177_ sky130_fd_sc_hd__mux2_1
XFILLER_109_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13150_ clknet_leaf_167_clk _01844_ VGND VGND VPWR VPWR tag_array.tag1\[8\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_10362_ net752 net3140 net539 VGND VGND VPWR VPWR _02109_ sky130_fd_sc_hd__mux2_1
XFILLER_3_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12101_ clknet_leaf_77_clk _00909_ VGND VGND VPWR VPWR data_array.data1\[14\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_151_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10293_ net1948 net991 net640 VGND VGND VPWR VPWR _02040_ sky130_fd_sc_hd__mux2_1
X_13081_ clknet_leaf_264_clk _01775_ VGND VGND VPWR VPWR data_array.data1\[13\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
X_12032_ clknet_leaf_92_clk _00840_ VGND VGND VPWR VPWR data_array.data0\[6\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold190 data_array.data0\[2\]\[20\] VGND VGND VPWR VPWR net1841 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_72_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1602 net1603 VGND VGND VPWR VPWR net1602 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_72_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1613 _03508_ VGND VGND VPWR VPWR net1613 sky130_fd_sc_hd__clkbuf_4
Xfanout1624 net1627 VGND VGND VPWR VPWR net1624 sky130_fd_sc_hd__buf_2
XFILLER_104_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1635 net1637 VGND VGND VPWR VPWR net1635 sky130_fd_sc_hd__clkbuf_4
Xfanout1646 net1647 VGND VGND VPWR VPWR net1646 sky130_fd_sc_hd__clkbuf_2
XFILLER_120_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout670 _05549_ VGND VGND VPWR VPWR net670 sky130_fd_sc_hd__clkbuf_4
Xfanout681 net685 VGND VGND VPWR VPWR net681 sky130_fd_sc_hd__clkbuf_8
XFILLER_77_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout692 _05417_ VGND VGND VPWR VPWR net692 sky130_fd_sc_hd__buf_4
X_13983_ clknet_leaf_204_clk _02612_ VGND VGND VPWR VPWR data_array.data1\[5\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_830 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12934_ clknet_leaf_73_clk _01628_ VGND VGND VPWR VPWR data_array.data0\[13\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12865_ clknet_leaf_72_clk _01559_ VGND VGND VPWR VPWR data_array.data0\[12\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11816_ clknet_leaf_48_clk _00624_ VGND VGND VPWR VPWR data_array.data0\[7\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_12796_ clknet_leaf_231_clk _01490_ VGND VGND VPWR VPWR tag_array.tag1\[10\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_155_3334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_3345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ clknet_leaf_192_clk _00555_ VGND VGND VPWR VPWR data_array.data0\[8\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_159_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14466_ clknet_leaf_246_clk _03089_ VGND VGND VPWR VPWR data_array.data1\[7\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_172_3670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11678_ clknet_leaf_100_clk _00486_ VGND VGND VPWR VPWR tag_array.tag1\[1\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_116_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13417_ clknet_leaf_213_clk _02047_ VGND VGND VPWR VPWR data_array.data1\[8\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
X_10629_ net2074 net944 net466 VGND VGND VPWR VPWR _02374_ sky130_fd_sc_hd__mux2_1
X_14397_ clknet_leaf_79_clk _03020_ VGND VGND VPWR VPWR data_array.data1\[10\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13348_ clknet_leaf_230_clk _01978_ VGND VGND VPWR VPWR data_array.data0\[10\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
Xmax_cap826 _03347_ VGND VGND VPWR VPWR net826 sky130_fd_sc_hd__buf_1
XFILLER_170_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13279_ clknet_leaf_223_clk _01909_ VGND VGND VPWR VPWR data_array.data0\[11\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_130_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2508 tag_array.dirty0\[4\] VGND VGND VPWR VPWR net4159 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2519 tag_array.tag1\[12\]\[20\] VGND VGND VPWR VPWR net4170 sky130_fd_sc_hd__dlygate4sd3_1
X_07840_ data_array.data1\[4\]\[36\] net1414 net1320 data_array.data1\[7\]\[36\] _05044_
+ VGND VGND VPWR VPWR _05045_ sky130_fd_sc_hd__a221o_1
Xhold1807 data_array.data1\[15\]\[10\] VGND VGND VPWR VPWR net3458 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1818 data_array.data0\[10\]\[57\] VGND VGND VPWR VPWR net3469 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_679 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1829 tag_array.tag0\[3\]\[8\] VGND VGND VPWR VPWR net3480 sky130_fd_sc_hd__dlygate4sd3_1
X_07771_ data_array.data1\[9\]\[30\] net1583 net1487 data_array.data1\[10\]\[30\]
+ VGND VGND VPWR VPWR _04982_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_179_3802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09510_ net790 net2375 net621 VGND VGND VPWR VPWR _01263_ sky130_fd_sc_hd__mux2_1
X_06722_ tag_array.tag1\[0\]\[23\] net1419 net1325 tag_array.tag1\[3\]\[23\] _04028_
+ VGND VGND VPWR VPWR _04029_ sky130_fd_sc_hd__a221o_1
XFILLER_52_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09441_ net900 net3852 net582 VGND VGND VPWR VPWR _01194_ sky130_fd_sc_hd__mux2_1
X_06653_ tag_array.tag1\[9\]\[17\] net1607 net1511 tag_array.tag1\[10\]\[17\] VGND
+ VGND VPWR VPWR _03966_ sky130_fd_sc_hd__a22o_1
XFILLER_64_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09372_ net912 net2489 net407 VGND VGND VPWR VPWR _01125_ sky130_fd_sc_hd__mux2_1
X_06584_ tag_array.tag1\[8\]\[11\] net1388 net1294 tag_array.tag1\[11\]\[11\] _03902_
+ VGND VGND VPWR VPWR _03903_ sky130_fd_sc_hd__a221o_1
XFILLER_80_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08323_ net1125 _05451_ VGND VGND VPWR VPWR _05452_ sky130_fd_sc_hd__and2_1
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08254_ _03143_ _03147_ VGND VGND VPWR VPWR _05404_ sky130_fd_sc_hd__nor2_1
XFILLER_166_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07205_ data_array.data0\[1\]\[42\] net1579 net1483 data_array.data0\[2\]\[42\] VGND
+ VGND VPWR VPWR _04468_ sky130_fd_sc_hd__a22o_1
XFILLER_165_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08185_ fsm.state\[2\] net840 _05355_ VGND VGND VPWR VPWR _05356_ sky130_fd_sc_hd__a21o_1
XFILLER_4_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07136_ data_array.data0\[4\]\[36\] net1413 net1319 data_array.data0\[7\]\[36\] _04404_
+ VGND VGND VPWR VPWR _04405_ sky130_fd_sc_hd__a221o_1
XFILLER_174_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07067_ data_array.data0\[9\]\[30\] net1583 net1487 data_array.data0\[10\]\[30\]
+ VGND VGND VPWR VPWR _04342_ sky130_fd_sc_hd__a22o_1
Xoutput240 net240 VGND VGND VPWR VPWR mem_addr[19] sky130_fd_sc_hd__buf_2
Xoutput251 net251 VGND VGND VPWR VPWR mem_addr[29] sky130_fd_sc_hd__buf_2
X_06018_ data_array.rdata1\[62\] net1657 net843 VGND VGND VPWR VPWR _03473_ sky130_fd_sc_hd__a21o_1
XFILLER_0_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput262 net1164 VGND VGND VPWR VPWR mem_read sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput273 net273 VGND VGND VPWR VPWR mem_wdata[19] sky130_fd_sc_hd__buf_2
XFILLER_0_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput284 net284 VGND VGND VPWR VPWR mem_wdata[29] sky130_fd_sc_hd__buf_2
Xoutput295 net295 VGND VGND VPWR VPWR mem_wdata[39] sky130_fd_sc_hd__buf_2
XFILLER_58_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07969_ data_array.data1\[9\]\[48\] net1590 net1494 data_array.data1\[10\]\[48\]
+ VGND VGND VPWR VPWR _05162_ sky130_fd_sc_hd__a22o_1
XFILLER_74_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09708_ net754 net3574 net611 VGND VGND VPWR VPWR _01460_ sky130_fd_sc_hd__mux2_1
X_10980_ net3397 net1081 net343 VGND VGND VPWR VPWR _02724_ sky130_fd_sc_hd__mux2_1
XFILLER_74_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09639_ net733 net4289 net616 VGND VGND VPWR VPWR _01391_ sky130_fd_sc_hd__mux2_1
XFILLER_15_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12650_ clknet_leaf_261_clk _01344_ VGND VGND VPWR VPWR data_array.data0\[15\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11601_ clknet_leaf_128_clk _00409_ VGND VGND VPWR VPWR tag_array.tag1\[4\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12581_ clknet_leaf_138_clk _01275_ VGND VGND VPWR VPWR tag_array.tag0\[10\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14320_ clknet_leaf_122_clk _02949_ VGND VGND VPWR VPWR data_array.data1\[11\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11532_ clknet_leaf_172_clk _00340_ VGND VGND VPWR VPWR tag_array.valid1\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_156_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14251_ clknet_leaf_259_clk _02880_ VGND VGND VPWR VPWR data_array.data1\[12\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11463_ clknet_leaf_223_clk _00273_ VGND VGND VPWR VPWR data_array.data0\[0\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_150_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13202_ clknet_leaf_253_clk _00096_ VGND VGND VPWR VPWR data_array.rdata1\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10414_ net3171 net997 net663 VGND VGND VPWR VPWR _02160_ sky130_fd_sc_hd__mux2_1
X_14182_ clknet_leaf_59_clk _02811_ VGND VGND VPWR VPWR data_array.data0\[2\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_137_684 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11394_ clknet_leaf_139_clk _00204_ VGND VGND VPWR VPWR tag_array.tag1\[7\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_74_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13133_ clknet_leaf_168_clk _01827_ VGND VGND VPWR VPWR tag_array.tag0\[3\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_111_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10345_ net721 net3668 net594 VGND VGND VPWR VPWR _02092_ sky130_fd_sc_hd__mux2_1
XFILLER_151_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13064_ clknet_leaf_70_clk _01758_ VGND VGND VPWR VPWR data_array.data1\[13\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_10276_ net2066 net1057 net637 VGND VGND VPWR VPWR _02023_ sky130_fd_sc_hd__mux2_1
XFILLER_3_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12015_ clknet_leaf_270_clk _00823_ VGND VGND VPWR VPWR data_array.data0\[6\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout1410 net1422 VGND VGND VPWR VPWR net1410 sky130_fd_sc_hd__buf_2
Xfanout1421 net1422 VGND VGND VPWR VPWR net1421 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_5_11__f_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_5_11__leaf_clk sky130_fd_sc_hd__clkbuf_16
Xfanout1432 net1433 VGND VGND VPWR VPWR net1432 sky130_fd_sc_hd__clkbuf_4
Xfanout1443 net1447 VGND VGND VPWR VPWR net1443 sky130_fd_sc_hd__clkbuf_2
Xfanout1454 net1455 VGND VGND VPWR VPWR net1454 sky130_fd_sc_hd__clkbuf_4
XFILLER_66_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1465 net1467 VGND VGND VPWR VPWR net1465 sky130_fd_sc_hd__clkbuf_4
Xfanout1476 net1477 VGND VGND VPWR VPWR net1476 sky130_fd_sc_hd__clkbuf_4
XFILLER_120_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1487 net1488 VGND VGND VPWR VPWR net1487 sky130_fd_sc_hd__clkbuf_4
Xfanout1498 net1517 VGND VGND VPWR VPWR net1498 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_109_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_543 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13966_ clknet_leaf_269_clk _02595_ VGND VGND VPWR VPWR data_array.data1\[5\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_126_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12917_ clknet_leaf_226_clk _01611_ VGND VGND VPWR VPWR data_array.data0\[13\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13897_ clknet_leaf_266_clk _02526_ VGND VGND VPWR VPWR data_array.data1\[4\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_94_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_100_Left_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12848_ clknet_leaf_222_clk _01542_ VGND VGND VPWR VPWR data_array.data0\[12\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12779_ clknet_leaf_178_clk _01473_ VGND VGND VPWR VPWR tag_array.tag0\[6\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_170_3629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_746 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14449_ clknet_leaf_73_clk _03072_ VGND VGND VPWR VPWR data_array.data1\[7\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold904 data_array.data0\[1\]\[35\] VGND VGND VPWR VPWR net2555 sky130_fd_sc_hd__dlygate4sd3_1
Xhold915 data_array.data0\[4\]\[47\] VGND VGND VPWR VPWR net2566 sky130_fd_sc_hd__dlygate4sd3_1
Xhold926 data_array.data1\[2\]\[7\] VGND VGND VPWR VPWR net2577 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold937 tag_array.tag0\[13\]\[22\] VGND VGND VPWR VPWR net2588 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold948 data_array.data1\[9\]\[55\] VGND VGND VPWR VPWR net2599 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_127_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09990_ net868 net3942 net377 VGND VGND VPWR VPWR _01739_ sky130_fd_sc_hd__mux2_1
Xhold959 tag_array.tag0\[14\]\[23\] VGND VGND VPWR VPWR net2610 sky130_fd_sc_hd__dlygate4sd3_1
X_08941_ net1003 net4363 net428 VGND VGND VPWR VPWR _00697_ sky130_fd_sc_hd__mux2_1
XFILLER_143_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2305 tag_array.tag0\[4\]\[18\] VGND VGND VPWR VPWR net3956 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_142_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2316 data_array.data0\[10\]\[43\] VGND VGND VPWR VPWR net3967 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08872_ net1018 net3641 net437 VGND VGND VPWR VPWR _00629_ sky130_fd_sc_hd__mux2_1
Xhold2327 data_array.data1\[13\]\[9\] VGND VGND VPWR VPWR net3978 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2338 data_array.data1\[13\]\[47\] VGND VGND VPWR VPWR net3989 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1604 tag_array.tag0\[14\]\[20\] VGND VGND VPWR VPWR net3255 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2349 tag_array.tag0\[11\]\[10\] VGND VGND VPWR VPWR net4000 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1615 data_array.data1\[15\]\[36\] VGND VGND VPWR VPWR net3266 sky130_fd_sc_hd__dlygate4sd3_1
X_07823_ net1189 _05023_ _05027_ net1615 VGND VGND VPWR VPWR _05030_ sky130_fd_sc_hd__a22o_1
XFILLER_97_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1626 tag_array.tag0\[1\]\[0\] VGND VGND VPWR VPWR net3277 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1637 tag_array.tag0\[5\]\[20\] VGND VGND VPWR VPWR net3288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1648 data_array.data1\[12\]\[48\] VGND VGND VPWR VPWR net3299 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1659 data_array.data1\[6\]\[20\] VGND VGND VPWR VPWR net3310 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07754_ data_array.data1\[12\]\[28\] net1349 net1255 data_array.data1\[15\]\[28\]
+ _04966_ VGND VGND VPWR VPWR _04967_ sky130_fd_sc_hd__a221o_1
XFILLER_65_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06705_ tag_array.tag1\[12\]\[22\] net1362 net1268 tag_array.tag1\[15\]\[22\] _04012_
+ VGND VGND VPWR VPWR _04013_ sky130_fd_sc_hd__a221o_1
XFILLER_65_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07685_ data_array.data1\[1\]\[22\] net1537 net1441 data_array.data1\[2\]\[22\] VGND
+ VGND VPWR VPWR _04904_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_91_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_91_clk sky130_fd_sc_hd__clkbuf_8
X_09424_ net968 net3913 net578 VGND VGND VPWR VPWR _01177_ sky130_fd_sc_hd__mux2_1
X_06636_ net1229 _03945_ _03949_ net1187 VGND VGND VPWR VPWR _03951_ sky130_fd_sc_hd__a22o_1
X_09355_ net982 net3150 net402 VGND VGND VPWR VPWR _01108_ sky130_fd_sc_hd__mux2_1
X_06567_ tag_array.tag1\[1\]\[9\] net1607 net1511 tag_array.tag1\[2\]\[9\] VGND VGND
+ VPWR VPWR _03888_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_47_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08306_ net2320 net1068 net693 VGND VGND VPWR VPWR _00231_ sky130_fd_sc_hd__mux2_1
XFILLER_100_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09286_ net734 net4268 net557 VGND VGND VPWR VPWR _01040_ sky130_fd_sc_hd__mux2_1
XFILLER_139_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06498_ tag_array.tag1\[4\]\[3\] net1371 net1277 tag_array.tag1\[7\]\[3\] _03824_
+ VGND VGND VPWR VPWR _03825_ sky130_fd_sc_hd__a221o_1
XFILLER_165_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08237_ fsm.tag_out1\[14\] net816 net808 fsm.tag_out0\[14\] _05392_ VGND VGND VPWR
+ VPWR _05393_ sky130_fd_sc_hd__a221o_1
XFILLER_119_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08168_ lru_array.lru_mem\[12\] net1373 net1279 lru_array.lru_mem\[15\] _05342_ VGND
+ VGND VPWR VPWR _05343_ sky130_fd_sc_hd__a221o_1
XFILLER_106_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_91_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07119_ net1188 _04383_ _04387_ net1614 VGND VGND VPWR VPWR _04390_ sky130_fd_sc_hd__a22o_1
X_08099_ net1225 _05275_ _05279_ net1177 VGND VGND VPWR VPWR _05281_ sky130_fd_sc_hd__a22o_1
XFILLER_122_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10130_ net1026 net4055 net364 VGND VGND VPWR VPWR _01878_ sky130_fd_sc_hd__mux2_1
XFILLER_69_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10061_ net779 net3839 net599 VGND VGND VPWR VPWR _01810_ sky130_fd_sc_hd__mux2_1
XFILLER_0_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2850 data_array.data0\[9\]\[58\] VGND VGND VPWR VPWR net4501 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_125_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2861 tag_array.tag0\[7\]\[5\] VGND VGND VPWR VPWR net4512 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2872 data_array.data0\[14\]\[42\] VGND VGND VPWR VPWR net4523 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_47_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2883 tag_array.tag0\[9\]\[6\] VGND VGND VPWR VPWR net4534 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2894 data_array.data1\[11\]\[2\] VGND VGND VPWR VPWR net4545 sky130_fd_sc_hd__dlygate4sd3_1
X_13820_ clknet_leaf_212_clk _02449_ VGND VGND VPWR VPWR data_array.data1\[2\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13751_ clknet_leaf_78_clk _02380_ VGND VGND VPWR VPWR data_array.data1\[1\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
X_10963_ net890 net3433 net527 VGND VGND VPWR VPWR _02708_ sky130_fd_sc_hd__mux2_1
XFILLER_90_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_82_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_82_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_67_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12702_ clknet_leaf_170_clk _01396_ VGND VGND VPWR VPWR tag_array.tag0\[8\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_67_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13682_ clknet_leaf_84_clk _02311_ VGND VGND VPWR VPWR data_array.data1\[15\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_44_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10894_ net908 net2756 net514 VGND VGND VPWR VPWR _02639_ sky130_fd_sc_hd__mux2_1
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12633_ clknet_leaf_63_clk _01327_ VGND VGND VPWR VPWR data_array.data0\[15\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_84_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12564_ clknet_leaf_155_clk _01258_ VGND VGND VPWR VPWR tag_array.tag0\[11\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_180_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14303_ clknet_leaf_194_clk _02932_ VGND VGND VPWR VPWR data_array.data1\[11\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11515_ clknet_leaf_231_clk _00323_ VGND VGND VPWR VPWR tag_array.tag1\[9\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_12495_ clknet_leaf_79_clk _01189_ VGND VGND VPWR VPWR data_array.data1\[9\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_157_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14234_ clknet_leaf_46_clk _02863_ VGND VGND VPWR VPWR data_array.data1\[12\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_156_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11446_ clknet_leaf_245_clk _00256_ VGND VGND VPWR VPWR data_array.data0\[0\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14165_ clknet_leaf_225_clk _02794_ VGND VGND VPWR VPWR data_array.data0\[2\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11377_ net820 net3440 _05562_ VGND VGND VPWR VPWR _03120_ sky130_fd_sc_hd__mux2_1
XFILLER_98_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13116_ clknet_leaf_177_clk _01810_ VGND VGND VPWR VPWR tag_array.tag0\[3\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_10328_ net788 net4455 net591 VGND VGND VPWR VPWR _02075_ sky130_fd_sc_hd__mux2_1
X_14096_ clknet_leaf_14_clk _02725_ VGND VGND VPWR VPWR data_array.data0\[1\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_140_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_167_3580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ clknet_leaf_110_clk _01741_ VGND VGND VPWR VPWR data_array.data0\[3\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
X_10259_ net708 net1922 net596 VGND VGND VPWR VPWR _02006_ sky130_fd_sc_hd__mux2_1
XFILLER_61_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1240 net1282 VGND VGND VPWR VPWR net1240 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_128_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1251 net1258 VGND VGND VPWR VPWR net1251 sky130_fd_sc_hd__clkbuf_4
Xfanout1262 net1264 VGND VGND VPWR VPWR net1262 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_163_3488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1273 net1282 VGND VGND VPWR VPWR net1273 sky130_fd_sc_hd__clkbuf_2
XFILLER_94_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_163_3499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1284 net1289 VGND VGND VPWR VPWR net1284 sky130_fd_sc_hd__clkbuf_4
Xfanout1295 net1298 VGND VGND VPWR VPWR net1295 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_124_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13949_ clknet_leaf_5_clk _02578_ VGND VGND VPWR VPWR data_array.data1\[4\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_73_clk clknet_5_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_73_clk sky130_fd_sc_hd__clkbuf_8
X_07470_ data_array.data1\[0\]\[2\] net1336 net1242 data_array.data1\[3\]\[2\] _04708_
+ VGND VGND VPWR VPWR _04709_ sky130_fd_sc_hd__a221o_1
X_06421_ tag_array.tag0\[4\]\[21\] net1407 net1313 tag_array.tag0\[7\]\[21\] _03754_
+ VGND VGND VPWR VPWR _03755_ sky130_fd_sc_hd__a221o_1
XFILLER_34_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09140_ net981 net4212 net566 VGND VGND VPWR VPWR _00894_ sky130_fd_sc_hd__mux2_1
X_06352_ tag_array.tag0\[13\]\[15\] net1593 net1497 tag_array.tag0\[14\]\[15\] VGND
+ VGND VPWR VPWR _03692_ sky130_fd_sc_hd__a22o_1
XFILLER_175_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09071_ net1003 net4424 net412 VGND VGND VPWR VPWR _00825_ sky130_fd_sc_hd__mux2_1
X_06283_ net1634 _03623_ _03627_ net1208 VGND VGND VPWR VPWR _03630_ sky130_fd_sc_hd__a22o_1
XFILLER_30_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08022_ net1170 _05205_ _05209_ net1218 VGND VGND VPWR VPWR _05211_ sky130_fd_sc_hd__a22o_1
XFILLER_163_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold701 data_array.data1\[13\]\[44\] VGND VGND VPWR VPWR net2352 sky130_fd_sc_hd__dlygate4sd3_1
Xhold712 data_array.data1\[4\]\[3\] VGND VGND VPWR VPWR net2363 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold723 tag_array.tag0\[7\]\[13\] VGND VGND VPWR VPWR net2374 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_157_1031 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold734 data_array.data1\[1\]\[39\] VGND VGND VPWR VPWR net2385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold745 data_array.data1\[5\]\[10\] VGND VGND VPWR VPWR net2396 sky130_fd_sc_hd__dlygate4sd3_1
Xhold756 data_array.data0\[7\]\[37\] VGND VGND VPWR VPWR net2407 sky130_fd_sc_hd__dlygate4sd3_1
Xhold767 data_array.data0\[0\]\[38\] VGND VGND VPWR VPWR net2418 sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 data_array.data0\[1\]\[43\] VGND VGND VPWR VPWR net2429 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09973_ net936 net3400 net376 VGND VGND VPWR VPWR _01722_ sky130_fd_sc_hd__mux2_1
Xhold789 data_array.data0\[1\]\[10\] VGND VGND VPWR VPWR net2440 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2102 tag_array.tag0\[5\]\[7\] VGND VGND VPWR VPWR net3753 sky130_fd_sc_hd__dlygate4sd3_1
X_08924_ net1068 net2870 net432 VGND VGND VPWR VPWR _00680_ sky130_fd_sc_hd__mux2_1
Xhold2113 data_array.data1\[11\]\[27\] VGND VGND VPWR VPWR net3764 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2124 data_array.data1\[3\]\[44\] VGND VGND VPWR VPWR net3775 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2135 data_array.data0\[12\]\[21\] VGND VGND VPWR VPWR net3786 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1401 data_array.data0\[11\]\[46\] VGND VGND VPWR VPWR net3052 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2146 data_array.data0\[5\]\[13\] VGND VGND VPWR VPWR net3797 sky130_fd_sc_hd__dlygate4sd3_1
X_08855_ net1085 net4059 net434 VGND VGND VPWR VPWR _00612_ sky130_fd_sc_hd__mux2_1
Xhold2157 tag_array.tag0\[1\]\[4\] VGND VGND VPWR VPWR net3808 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1412 tag_array.tag1\[15\]\[1\] VGND VGND VPWR VPWR net3063 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1423 tag_array.dirty0\[11\] VGND VGND VPWR VPWR net3074 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2168 tag_array.dirty0\[9\] VGND VGND VPWR VPWR net3819 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1434 data_array.data1\[13\]\[12\] VGND VGND VPWR VPWR net3085 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2179 tag_array.tag0\[12\]\[21\] VGND VGND VPWR VPWR net3830 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1445 data_array.data1\[15\]\[55\] VGND VGND VPWR VPWR net3096 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07806_ data_array.data1\[1\]\[33\] net1587 net1491 data_array.data1\[2\]\[33\] VGND
+ VGND VPWR VPWR _05014_ sky130_fd_sc_hd__a22o_1
Xhold1456 data_array.data1\[14\]\[16\] VGND VGND VPWR VPWR net3107 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_88_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08786_ net2694 net1103 net444 VGND VGND VPWR VPWR _00544_ sky130_fd_sc_hd__mux2_1
Xhold1467 tag_array.tag0\[13\]\[9\] VGND VGND VPWR VPWR net3118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1478 data_array.data1\[12\]\[25\] VGND VGND VPWR VPWR net3129 sky130_fd_sc_hd__dlygate4sd3_1
X_05998_ net149 net1154 _03458_ _03459_ VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__a22o_1
XFILLER_26_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1489 tag_array.tag0\[15\]\[10\] VGND VGND VPWR VPWR net3140 sky130_fd_sc_hd__dlygate4sd3_1
X_07737_ _04950_ _04951_ VGND VGND VPWR VPWR _00082_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_49_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_64_clk clknet_5_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_64_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_81_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07668_ data_array.data1\[0\]\[20\] net1419 net1325 data_array.data1\[3\]\[20\] _04888_
+ VGND VGND VPWR VPWR _04889_ sky130_fd_sc_hd__a221o_1
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09407_ net1039 net2865 net580 VGND VGND VPWR VPWR _01160_ sky130_fd_sc_hd__mux2_1
XFILLER_41_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06619_ tag_array.tag1\[0\]\[14\] net1368 net1274 tag_array.tag1\[3\]\[14\] _03934_
+ VGND VGND VPWR VPWR _03935_ sky130_fd_sc_hd__a221o_1
XFILLER_13_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07599_ data_array.data1\[13\]\[14\] net1572 net1476 data_array.data1\[14\]\[14\]
+ VGND VGND VPWR VPWR _04826_ sky130_fd_sc_hd__a22o_1
X_09338_ net1049 net3452 net407 VGND VGND VPWR VPWR _01091_ sky130_fd_sc_hd__mux2_1
XFILLER_179_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09269_ net703 net2897 net570 VGND VGND VPWR VPWR _01023_ sky130_fd_sc_hd__mux2_1
XFILLER_126_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11300_ net1094 net3902 net801 VGND VGND VPWR VPWR _03043_ sky130_fd_sc_hd__mux2_1
XFILLER_181_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12280_ clknet_leaf_168_clk _01038_ VGND VGND VPWR VPWR tag_array.tag1\[13\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11231_ net1104 net3296 net673 VGND VGND VPWR VPWR _02974_ sky130_fd_sc_hd__mux2_1
XFILLER_106_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11162_ net871 net3163 net551 VGND VGND VPWR VPWR _02905_ sky130_fd_sc_hd__mux2_1
XFILLER_20_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10113_ net1093 net4429 net366 VGND VGND VPWR VPWR _01861_ sky130_fd_sc_hd__mux2_1
XFILLER_1_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11093_ net2353 net888 net329 VGND VGND VPWR VPWR _02836_ sky130_fd_sc_hd__mux2_1
X_10044_ net908 net2722 net555 VGND VGND VPWR VPWR _01793_ sky130_fd_sc_hd__mux2_1
XFILLER_96_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold50 tag_array.valid1\[11\] VGND VGND VPWR VPWR net1701 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2680 data_array.data1\[15\]\[40\] VGND VGND VPWR VPWR net4331 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_69_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold61 tag_array.valid0\[2\] VGND VGND VPWR VPWR net1712 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 tag_array.valid1\[1\] VGND VGND VPWR VPWR net1723 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_69_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold83 data_array.data0\[1\]\[19\] VGND VGND VPWR VPWR net1734 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2691 tag_array.tag1\[3\]\[2\] VGND VGND VPWR VPWR net4342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 tag_array.tag1\[2\]\[6\] VGND VGND VPWR VPWR net1745 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13803_ clknet_leaf_257_clk _02432_ VGND VGND VPWR VPWR data_array.data1\[2\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1990 data_array.data0\[7\]\[23\] VGND VGND VPWR VPWR net3641 sky130_fd_sc_hd__dlygate4sd3_1
X_11995_ clknet_leaf_209_clk _00803_ VGND VGND VPWR VPWR data_array.data0\[6\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_55_clk clknet_5_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_55_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_28_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13734_ clknet_leaf_70_clk _02363_ VGND VGND VPWR VPWR data_array.data1\[1\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_10946_ net958 net4174 net533 VGND VGND VPWR VPWR _02691_ sky130_fd_sc_hd__mux2_1
XFILLER_90_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13665_ clknet_leaf_263_clk _02294_ VGND VGND VPWR VPWR data_array.data1\[15\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_10877_ net978 net3586 net521 VGND VGND VPWR VPWR _02622_ sky130_fd_sc_hd__mux2_1
XFILLER_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12616_ clknet_leaf_127_clk _01310_ VGND VGND VPWR VPWR tag_array.tag0\[0\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_13596_ clknet_leaf_228_clk _02225_ VGND VGND VPWR VPWR data_array.data0\[9\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_12547_ clknet_leaf_178_clk _01241_ VGND VGND VPWR VPWR tag_array.tag0\[11\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_145_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12478_ clknet_leaf_67_clk _01172_ VGND VGND VPWR VPWR data_array.data1\[9\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_3 _00078_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14217_ clknet_leaf_264_clk _02846_ VGND VGND VPWR VPWR data_array.data1\[12\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11429_ clknet_leaf_15_clk _00239_ VGND VGND VPWR VPWR data_array.data0\[0\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_5_9__f_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_5_9__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_125_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14148_ clknet_leaf_114_clk _02777_ VGND VGND VPWR VPWR data_array.data0\[1\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_165_3528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_165_3539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06970_ data_array.data0\[1\]\[21\] net1556 net1460 data_array.data0\[2\]\[21\] VGND
+ VGND VPWR VPWR _04254_ sky130_fd_sc_hd__a22o_1
X_14079_ clknet_leaf_17_clk _02708_ VGND VGND VPWR VPWR data_array.data1\[6\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_101_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_182_3853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_3864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05921_ data_array.rdata0\[30\] net850 net1147 VGND VGND VPWR VPWR _03408_ sky130_fd_sc_hd__o21a_1
XFILLER_6_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1070 net1071 VGND VGND VPWR VPWR net1070 sky130_fd_sc_hd__clkbuf_2
X_08640_ net2306 net764 net510 VGND VGND VPWR VPWR _00399_ sky130_fd_sc_hd__mux2_1
Xfanout1081 _05434_ VGND VGND VPWR VPWR net1081 sky130_fd_sc_hd__dlymetal6s2s_1
X_05852_ data_array.rdata0\[7\] net1659 net1149 VGND VGND VPWR VPWR _03362_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_175_Right_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1092 net1093 VGND VGND VPWR VPWR net1092 sky130_fd_sc_hd__clkbuf_2
XFILLER_81_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_736 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08571_ net1713 net506 VGND VGND VPWR VPWR _00336_ sky130_fd_sc_hd__or2_1
X_05783_ net10 fsm.tag_out1\[11\] VGND VGND VPWR VPWR _03300_ sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_46_clk clknet_5_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_46_clk sky130_fd_sc_hd__clkbuf_8
X_07522_ data_array.data1\[13\]\[7\] net1589 net1493 data_array.data1\[14\]\[7\] VGND
+ VGND VPWR VPWR _04756_ sky130_fd_sc_hd__a22o_1
XFILLER_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07453_ data_array.data1\[12\]\[1\] net1330 net1236 data_array.data1\[15\]\[1\] _04692_
+ VGND VGND VPWR VPWR _04693_ sky130_fd_sc_hd__a221o_1
XFILLER_37_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06404_ net1208 _03733_ _03737_ net1634 VGND VGND VPWR VPWR _03740_ sky130_fd_sc_hd__a22o_1
X_07384_ net1170 _04625_ _04629_ net1218 VGND VGND VPWR VPWR _04631_ sky130_fd_sc_hd__a22o_1
XFILLER_163_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09123_ net1050 net2720 net574 VGND VGND VPWR VPWR _00877_ sky130_fd_sc_hd__mux2_1
X_06335_ tag_array.tag0\[12\]\[13\] net1410 net1316 tag_array.tag0\[15\]\[13\] _03676_
+ VGND VGND VPWR VPWR _03677_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_40_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09054_ net1068 net4001 net416 VGND VGND VPWR VPWR _00808_ sky130_fd_sc_hd__mux2_1
X_06266_ tag_array.tag0\[1\]\[7\] net1607 net1511 tag_array.tag0\[2\]\[7\] VGND VGND
+ VPWR VPWR _03614_ sky130_fd_sc_hd__a22o_1
X_08005_ data_array.data1\[4\]\[51\] net1334 net1240 data_array.data1\[7\]\[51\] _05194_
+ VGND VGND VPWR VPWR _05195_ sky130_fd_sc_hd__a221o_1
Xhold520 data_array.data0\[2\]\[12\] VGND VGND VPWR VPWR net2171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold531 tag_array.tag1\[2\]\[10\] VGND VGND VPWR VPWR net2182 sky130_fd_sc_hd__dlygate4sd3_1
X_06197_ _03550_ _03551_ VGND VGND VPWR VPWR _00131_ sky130_fd_sc_hd__or2_1
Xhold542 data_array.data0\[6\]\[2\] VGND VGND VPWR VPWR net2193 sky130_fd_sc_hd__dlygate4sd3_1
Xhold553 data_array.data0\[6\]\[26\] VGND VGND VPWR VPWR net2204 sky130_fd_sc_hd__dlygate4sd3_1
Xhold564 data_array.data1\[14\]\[62\] VGND VGND VPWR VPWR net2215 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold575 data_array.data0\[0\]\[35\] VGND VGND VPWR VPWR net2226 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold586 tag_array.tag1\[4\]\[4\] VGND VGND VPWR VPWR net2237 sky130_fd_sc_hd__dlygate4sd3_1
Xhold597 tag_array.tag1\[0\]\[4\] VGND VGND VPWR VPWR net2248 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09956_ net1007 net3647 net373 VGND VGND VPWR VPWR _01705_ sky130_fd_sc_hd__mux2_1
XFILLER_98_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08907_ net876 net2930 net437 VGND VGND VPWR VPWR _00664_ sky130_fd_sc_hd__mux2_1
XFILLER_66_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09887_ net920 net4388 net382 VGND VGND VPWR VPWR _01637_ sky130_fd_sc_hd__mux2_1
Xhold1220 tag_array.tag1\[0\]\[17\] VGND VGND VPWR VPWR net2871 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1231 data_array.data0\[10\]\[19\] VGND VGND VPWR VPWR net2882 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_86_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1242 data_array.data0\[12\]\[44\] VGND VGND VPWR VPWR net2893 sky130_fd_sc_hd__dlygate4sd3_1
X_08838_ net3146 net894 net444 VGND VGND VPWR VPWR _00596_ sky130_fd_sc_hd__mux2_1
Xhold1253 data_array.data0\[2\]\[45\] VGND VGND VPWR VPWR net2904 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_142_Right_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1264 tag_array.tag1\[5\]\[8\] VGND VGND VPWR VPWR net2915 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1275 tag_array.tag0\[6\]\[14\] VGND VGND VPWR VPWR net2926 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1286 tag_array.tag0\[14\]\[5\] VGND VGND VPWR VPWR net2937 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08769_ net749 net3627 net451 VGND VGND VPWR VPWR _00528_ sky130_fd_sc_hd__mux2_1
Xhold1297 data_array.data0\[14\]\[7\] VGND VGND VPWR VPWR net2948 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_140_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_37_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_8
X_10800_ net3176 net1030 net511 VGND VGND VPWR VPWR _02545_ sky130_fd_sc_hd__mux2_1
XFILLER_60_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11780_ clknet_leaf_23_clk _00588_ VGND VGND VPWR VPWR data_array.data0\[8\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_64_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10731_ net1050 net2595 net497 VGND VGND VPWR VPWR _02476_ sky130_fd_sc_hd__mux2_1
XFILLER_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13450_ clknet_leaf_179_clk _02080_ VGND VGND VPWR VPWR tag_array.tag0\[1\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_10662_ net1746 net1070 net487 VGND VGND VPWR VPWR _02407_ sky130_fd_sc_hd__mux2_1
XFILLER_167_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12401_ clknet_leaf_60_clk _01095_ VGND VGND VPWR VPWR data_array.data0\[14\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_13381_ clknet_leaf_265_clk _02011_ VGND VGND VPWR VPWR data_array.data1\[8\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_10593_ net1776 net1090 net470 VGND VGND VPWR VPWR _02338_ sky130_fd_sc_hd__mux2_1
XFILLER_139_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12332_ clknet_leaf_52_clk _00005_ VGND VGND VPWR VPWR data_array.rdata0\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_749 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12263_ clknet_leaf_234_clk _01021_ VGND VGND VPWR VPWR tag_array.tag1\[14\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_79_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14002_ clknet_leaf_87_clk _02631_ VGND VGND VPWR VPWR data_array.data1\[5\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
X_11214_ net919 net4519 net656 VGND VGND VPWR VPWR _02957_ sky130_fd_sc_hd__mux2_1
X_12194_ clknet_leaf_151_clk _00142_ VGND VGND VPWR VPWR fsm.tag_out0\[1\] sky130_fd_sc_hd__dfxtp_1
X_11145_ net938 net3892 net548 VGND VGND VPWR VPWR _02888_ sky130_fd_sc_hd__mux2_1
XFILLER_0_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11076_ net2751 net956 net333 VGND VGND VPWR VPWR _02819_ sky130_fd_sc_hd__mux2_1
Xinput140 mem_rdata[47] VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput151 mem_rdata[57] VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_1
X_10027_ net978 net3929 net562 VGND VGND VPWR VPWR _01776_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_160_3436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput162 mem_rdata[9] VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_160_3447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_28_clk clknet_5_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_8
X_11978_ clknet_leaf_208_clk _00786_ VGND VGND VPWR VPWR data_array.data0\[4\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13717_ clknet_leaf_200_clk _02346_ VGND VGND VPWR VPWR data_array.data1\[1\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_10929_ net1024 net4561 net529 VGND VGND VPWR VPWR _02674_ sky130_fd_sc_hd__mux2_1
XFILLER_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13648_ clknet_leaf_19_clk _02277_ VGND VGND VPWR VPWR data_array.data1\[15\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_119_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13579_ clknet_leaf_73_clk _02208_ VGND VGND VPWR VPWR data_array.data0\[9\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_158_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06120_ data_array.rdata0\[35\] net1135 net1113 data_array.rdata1\[35\] VGND VGND
+ VPWR VPWR net291 sky130_fd_sc_hd__a22o_1
XFILLER_8_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06051_ net1162 net7 fsm.tag_out1\[8\] net1132 VGND VGND VPWR VPWR _03489_ sky130_fd_sc_hd__a22o_1
XFILLER_172_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_184_3904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_184_3915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_99_Right_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09810_ net970 net2631 net387 VGND VGND VPWR VPWR _01561_ sky130_fd_sc_hd__mux2_1
XFILLER_67_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout329 net332 VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__buf_4
XFILLER_113_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1078 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09741_ net724 net3272 net683 VGND VGND VPWR VPWR _01493_ sky130_fd_sc_hd__mux2_1
X_06953_ data_array.data0\[0\]\[19\] net1389 net1295 data_array.data0\[3\]\[19\] _04238_
+ VGND VGND VPWR VPWR _04239_ sky130_fd_sc_hd__a221o_1
X_05904_ data_array.rdata1\[24\] net832 net841 VGND VGND VPWR VPWR _03397_ sky130_fd_sc_hd__a21o_1
X_09672_ net698 net2533 net613 VGND VGND VPWR VPWR _01424_ sky130_fd_sc_hd__mux2_1
X_06884_ data_array.data0\[9\]\[13\] net1553 net1457 data_array.data0\[10\]\[13\]
+ VGND VGND VPWR VPWR _04176_ sky130_fd_sc_hd__a22o_1
XFILLER_82_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08623_ net730 net4425 net522 VGND VGND VPWR VPWR _00382_ sky130_fd_sc_hd__mux2_1
X_05835_ data_array.rdata1\[1\] net828 net837 VGND VGND VPWR VPWR _03351_ sky130_fd_sc_hd__a21o_1
XFILLER_54_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_19_clk clknet_5_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_8
X_08554_ net740 net3213 net589 VGND VGND VPWR VPWR _00322_ sky130_fd_sc_hd__mux2_1
X_05766_ net16 fsm.tag_out1\[16\] VGND VGND VPWR VPWR _03283_ sky130_fd_sc_hd__xor2_2
X_07505_ net1219 _04735_ _04739_ net1171 VGND VGND VPWR VPWR _04741_ sky130_fd_sc_hd__a22o_1
XFILLER_51_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08485_ net1705 net632 VGND VGND VPWR VPWR _00290_ sky130_fd_sc_hd__nand2b_1
X_05697_ _03167_ _03193_ VGND VGND VPWR VPWR _03214_ sky130_fd_sc_hd__or2_1
X_07436_ data_array.data0\[1\]\[63\] net1548 net1452 data_array.data0\[2\]\[63\] VGND
+ VGND VPWR VPWR _04678_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_21_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07367_ data_array.data0\[0\]\[57\] net1348 net1254 data_array.data0\[3\]\[57\] _04614_
+ VGND VGND VPWR VPWR _04615_ sky130_fd_sc_hd__a221o_1
XFILLER_164_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09106_ net860 net2302 net416 VGND VGND VPWR VPWR _00860_ sky130_fd_sc_hd__mux2_1
X_06318_ _03660_ _03661_ VGND VGND VPWR VPWR _00133_ sky130_fd_sc_hd__or2_1
XFILLER_176_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07298_ data_array.data0\[13\]\[51\] net1522 net1426 data_array.data0\[14\]\[51\]
+ VGND VGND VPWR VPWR _04552_ sky130_fd_sc_hd__a22o_1
XFILLER_175_192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09037_ net2624 net876 net421 VGND VGND VPWR VPWR _00792_ sky130_fd_sc_hd__mux2_1
XFILLER_124_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06249_ tag_array.tag0\[0\]\[5\] net1418 net1324 tag_array.tag0\[3\]\[5\] _03598_
+ VGND VGND VPWR VPWR _03599_ sky130_fd_sc_hd__a221o_1
XFILLER_151_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold350 data_array.data0\[8\]\[32\] VGND VGND VPWR VPWR net2001 sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 data_array.data1\[0\]\[3\] VGND VGND VPWR VPWR net2012 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold372 tag_array.tag1\[2\]\[15\] VGND VGND VPWR VPWR net2023 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold383 data_array.data0\[0\]\[42\] VGND VGND VPWR VPWR net2034 sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 data_array.data1\[1\]\[47\] VGND VGND VPWR VPWR net2045 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout830 net831 VGND VGND VPWR VPWR net830 sky130_fd_sc_hd__buf_6
XFILLER_131_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout841 net842 VGND VGND VPWR VPWR net841 sky130_fd_sc_hd__buf_6
Xfanout852 net853 VGND VGND VPWR VPWR net852 sky130_fd_sc_hd__buf_12
X_09939_ net1072 net3650 net375 VGND VGND VPWR VPWR _01688_ sky130_fd_sc_hd__mux2_1
Xfanout863 _05544_ VGND VGND VPWR VPWR net863 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_142_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout874 net875 VGND VGND VPWR VPWR net874 sky130_fd_sc_hd__clkbuf_2
Xfanout885 _05532_ VGND VGND VPWR VPWR net885 sky130_fd_sc_hd__buf_1
Xclkbuf_4_13_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_13_0_clk sky130_fd_sc_hd__clkbuf_8
X_12950_ clknet_leaf_220_clk _01644_ VGND VGND VPWR VPWR data_array.data0\[13\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout896 _05526_ VGND VGND VPWR VPWR net896 sky130_fd_sc_hd__clkbuf_2
Xhold1050 data_array.data0\[12\]\[9\] VGND VGND VPWR VPWR net2701 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1061 data_array.data1\[13\]\[7\] VGND VGND VPWR VPWR net2712 sky130_fd_sc_hd__dlygate4sd3_1
X_11901_ clknet_leaf_241_clk _00709_ VGND VGND VPWR VPWR data_array.data0\[5\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1072 data_array.data0\[11\]\[52\] VGND VGND VPWR VPWR net2723 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1083 data_array.data0\[9\]\[26\] VGND VGND VPWR VPWR net2734 sky130_fd_sc_hd__dlygate4sd3_1
X_12881_ clknet_leaf_54_clk _01575_ VGND VGND VPWR VPWR data_array.data0\[12\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_29_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1094 data_array.data1\[12\]\[45\] VGND VGND VPWR VPWR net2745 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11832_ clknet_leaf_11_clk _00640_ VGND VGND VPWR VPWR data_array.data0\[7\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11763_ clknet_leaf_54_clk _00571_ VGND VGND VPWR VPWR data_array.data0\[8\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10714_ net1799 net862 net487 VGND VGND VPWR VPWR _02459_ sky130_fd_sc_hd__mux2_1
X_13502_ clknet_leaf_35_clk _02131_ VGND VGND VPWR VPWR tag_array.dirty1\[8\] sky130_fd_sc_hd__dfxtp_1
X_14482_ clknet_leaf_165_clk _03105_ VGND VGND VPWR VPWR tag_array.dirty0\[1\] sky130_fd_sc_hd__dfxtp_1
X_11694_ clknet_leaf_105_clk _00502_ VGND VGND VPWR VPWR tag_array.tag1\[15\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_13433_ clknet_leaf_6_clk _02063_ VGND VGND VPWR VPWR data_array.data1\[8\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
X_10645_ net2059 net883 net466 VGND VGND VPWR VPWR _02390_ sky130_fd_sc_hd__mux2_1
Xclkload209 clknet_leaf_116_clk VGND VGND VPWR VPWR clkload209/Y sky130_fd_sc_hd__inv_6
X_13364_ clknet_leaf_160_clk _01994_ VGND VGND VPWR VPWR tag_array.tag0\[2\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_177_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10576_ net901 net3038 net457 VGND VGND VPWR VPWR _02321_ sky130_fd_sc_hd__mux2_1
X_12315_ clknet_leaf_196_clk _01073_ VGND VGND VPWR VPWR tag_array.tag1\[12\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_177_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13295_ clknet_leaf_73_clk _01925_ VGND VGND VPWR VPWR data_array.data0\[10\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_114_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12246_ clknet_leaf_191_clk _01004_ VGND VGND VPWR VPWR tag_array.tag1\[14\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_177_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12177_ clknet_leaf_158_clk _00985_ VGND VGND VPWR VPWR tag_array.tag0\[14\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_69_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11128_ net1004 net3178 net542 VGND VGND VPWR VPWR _02871_ sky130_fd_sc_hd__mux2_1
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11059_ net1783 net1027 net331 VGND VGND VPWR VPWR _02802_ sky130_fd_sc_hd__mux2_1
XFILLER_77_883 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1019 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_05620_ net18 VGND VGND VPWR VPWR _03142_ sky130_fd_sc_hd__inv_2
XFILLER_17_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_177_3752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_177_3763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_986 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08270_ fsm.state\[2\] net1644 net840 _05355_ VGND VGND VPWR VPWR _05415_ sky130_fd_sc_hd__a31o_1
XFILLER_32_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07221_ data_array.data0\[9\]\[44\] net1589 net1493 data_array.data0\[10\]\[44\]
+ VGND VGND VPWR VPWR _04482_ sky130_fd_sc_hd__a22o_1
XFILLER_34_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07152_ net1621 _04413_ _04417_ net1195 VGND VGND VPWR VPWR _04420_ sky130_fd_sc_hd__a22o_1
X_06103_ data_array.rdata0\[18\] net1135 net1112 data_array.rdata1\[18\] VGND VGND
+ VPWR VPWR net272 sky130_fd_sc_hd__a22o_1
XFILLER_121_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07083_ data_array.data0\[8\]\[31\] net1385 net1291 data_array.data0\[11\]\[31\]
+ _04356_ VGND VGND VPWR VPWR _04357_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_8_clk clknet_5_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_8
X_06034_ net1158 net1141 net1119 net29 VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__o31a_1
XFILLER_133_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07985_ data_array.data1\[8\]\[49\] net1382 net1288 data_array.data1\[11\]\[49\]
+ _05176_ VGND VGND VPWR VPWR _05177_ sky130_fd_sc_hd__a221o_1
XFILLER_101_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09724_ net791 net3254 net680 VGND VGND VPWR VPWR _01476_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06936_ data_array.data0\[8\]\[18\] net1377 net1283 data_array.data0\[11\]\[18\]
+ _04222_ VGND VGND VPWR VPWR _04223_ sky130_fd_sc_hd__a221o_1
XFILLER_170_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09655_ net769 net3825 net612 VGND VGND VPWR VPWR _01407_ sky130_fd_sc_hd__mux2_1
X_06867_ net1224 _04155_ _04159_ net1176 VGND VGND VPWR VPWR _04161_ sky130_fd_sc_hd__a22o_1
XFILLER_16_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08606_ net701 net3702 net536 VGND VGND VPWR VPWR _00365_ sky130_fd_sc_hd__mux2_1
XFILLER_27_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05818_ _03248_ _03265_ _03273_ _03278_ VGND VGND VPWR VPWR _03335_ sky130_fd_sc_hd__or4_1
X_09586_ net1006 net3127 net394 VGND VGND VPWR VPWR _01338_ sky130_fd_sc_hd__mux2_1
XFILLER_83_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06798_ data_array.data0\[5\]\[5\] net1545 net1449 data_array.data0\[6\]\[5\] VGND
+ VGND VPWR VPWR _04098_ sky130_fd_sc_hd__a22o_1
XFILLER_82_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08537_ net1279 net1200 VGND VGND VPWR VPWR _05595_ sky130_fd_sc_hd__nand2_1
XFILLER_179_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_05749_ net11 fsm.tag_out1\[12\] VGND VGND VPWR VPWR _03266_ sky130_fd_sc_hd__and2b_1
XFILLER_168_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08468_ net814 _05547_ net1699 VGND VGND VPWR VPWR _00285_ sky130_fd_sc_hd__a21o_1
XFILLER_144_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07419_ data_array.data0\[9\]\[62\] net1605 net1509 data_array.data0\[10\]\[62\]
+ VGND VGND VPWR VPWR _04662_ sky130_fd_sc_hd__a22o_1
X_08399_ net1991 net946 net686 VGND VGND VPWR VPWR _00262_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_98_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_682 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10430_ net1826 net934 net669 VGND VGND VPWR VPWR _02176_ sky130_fd_sc_hd__mux2_1
XFILLER_183_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10361_ net754 net2194 net539 VGND VGND VPWR VPWR _02108_ sky130_fd_sc_hd__mux2_1
XFILLER_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12100_ clknet_leaf_6_clk _00908_ VGND VGND VPWR VPWR data_array.data1\[14\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_76_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13080_ clknet_leaf_36_clk _01774_ VGND VGND VPWR VPWR data_array.data1\[13\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_163_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10292_ net2091 net994 net639 VGND VGND VPWR VPWR _02039_ sky130_fd_sc_hd__mux2_1
XFILLER_3_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12031_ clknet_leaf_244_clk _00839_ VGND VGND VPWR VPWR data_array.data0\[6\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold180 data_array.data1\[8\]\[52\] VGND VGND VPWR VPWR net1831 sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 data_array.data0\[8\]\[50\] VGND VGND VPWR VPWR net1842 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1603 net1612 VGND VGND VPWR VPWR net1603 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_72_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1614 net1617 VGND VGND VPWR VPWR net1614 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_72_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1625 net1627 VGND VGND VPWR VPWR net1625 sky130_fd_sc_hd__clkbuf_4
Xfanout1636 net1637 VGND VGND VPWR VPWR net1636 sky130_fd_sc_hd__buf_4
Xfanout1647 net1648 VGND VGND VPWR VPWR net1647 sky130_fd_sc_hd__buf_1
Xfanout660 _05551_ VGND VGND VPWR VPWR net660 sky130_fd_sc_hd__clkbuf_4
Xfanout671 net672 VGND VGND VPWR VPWR net671 sky130_fd_sc_hd__buf_4
XFILLER_144_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout682 net685 VGND VGND VPWR VPWR net682 sky130_fd_sc_hd__buf_2
Xfanout693 _05417_ VGND VGND VPWR VPWR net693 sky130_fd_sc_hd__buf_4
X_13982_ clknet_leaf_24_clk _02611_ VGND VGND VPWR VPWR data_array.data1\[5\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_842 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12933_ clknet_leaf_219_clk _01627_ VGND VGND VPWR VPWR data_array.data0\[13\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
X_12864_ clknet_leaf_260_clk _01558_ VGND VGND VPWR VPWR data_array.data0\[12\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_1030 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11815_ clknet_leaf_250_clk _00623_ VGND VGND VPWR VPWR data_array.data0\[7\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_12795_ clknet_leaf_134_clk _01489_ VGND VGND VPWR VPWR tag_array.tag1\[10\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_164_Left_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11746_ clknet_leaf_103_clk _00554_ VGND VGND VPWR VPWR data_array.data0\[8\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_155_3335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_155_3346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11677_ clknet_leaf_186_clk _00485_ VGND VGND VPWR VPWR tag_array.tag1\[1\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_14465_ clknet_leaf_55_clk _03088_ VGND VGND VPWR VPWR data_array.data1\[7\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_172_3660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13416_ clknet_leaf_118_clk _02046_ VGND VGND VPWR VPWR data_array.data1\[8\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
X_10628_ net2406 net950 net475 VGND VGND VPWR VPWR _02373_ sky130_fd_sc_hd__mux2_1
X_14396_ clknet_leaf_244_clk _03019_ VGND VGND VPWR VPWR data_array.data1\[10\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_133_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13347_ clknet_leaf_12_clk _01977_ VGND VGND VPWR VPWR data_array.data0\[10\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
X_10559_ net969 net4552 net453 VGND VGND VPWR VPWR _02304_ sky130_fd_sc_hd__mux2_1
XFILLER_115_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13278_ clknet_leaf_3_clk _01908_ VGND VGND VPWR VPWR data_array.data0\[11\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_173_Left_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12229_ clknet_leaf_151_clk _00158_ VGND VGND VPWR VPWR fsm.tag_out1\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_64_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2509 tag_array.tag1\[11\]\[1\] VGND VGND VPWR VPWR net4160 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1808 data_array.data0\[3\]\[23\] VGND VGND VPWR VPWR net3459 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1819 data_array.data1\[5\]\[55\] VGND VGND VPWR VPWR net3470 sky130_fd_sc_hd__dlygate4sd3_1
X_07770_ _04980_ _04981_ VGND VGND VPWR VPWR _00085_ sky130_fd_sc_hd__or2_1
X_06721_ tag_array.tag1\[1\]\[23\] net1610 net1514 tag_array.tag1\[2\]\[23\] VGND
+ VGND VPWR VPWR _04028_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_179_3803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09440_ net906 net4366 net578 VGND VGND VPWR VPWR _01193_ sky130_fd_sc_hd__mux2_1
X_06652_ tag_array.tag1\[4\]\[17\] net1418 net1324 tag_array.tag1\[7\]\[17\] _03964_
+ VGND VGND VPWR VPWR _03965_ sky130_fd_sc_hd__a221o_1
XFILLER_37_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_182_Left_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09371_ net916 net3950 net407 VGND VGND VPWR VPWR _01124_ sky130_fd_sc_hd__mux2_1
XFILLER_80_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06583_ tag_array.tag1\[9\]\[11\] net1575 net1479 tag_array.tag1\[10\]\[11\] VGND
+ VGND VPWR VPWR _03902_ sky130_fd_sc_hd__a22o_1
XFILLER_33_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08322_ net106 net41 net1643 VGND VGND VPWR VPWR _05451_ sky130_fd_sc_hd__mux2_1
XFILLER_178_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08253_ net714 net2316 net803 VGND VGND VPWR VPWR _00215_ sky130_fd_sc_hd__mux2_1
XFILLER_177_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07204_ data_array.data0\[12\]\[42\] net1395 net1301 data_array.data0\[15\]\[42\]
+ _04466_ VGND VGND VPWR VPWR _04467_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_31_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08184_ fsm.lru_out _03147_ VGND VGND VPWR VPWR _05355_ sky130_fd_sc_hd__nor2_1
XFILLER_181_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07135_ data_array.data0\[5\]\[36\] net1601 net1505 data_array.data0\[6\]\[36\] VGND
+ VGND VPWR VPWR _04404_ sky130_fd_sc_hd__a22o_1
XFILLER_118_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07066_ _04340_ _04341_ VGND VGND VPWR VPWR _00021_ sky130_fd_sc_hd__or2_1
Xoutput230 net230 VGND VGND VPWR VPWR mem_addr[0] sky130_fd_sc_hd__buf_2
XFILLER_134_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput241 net241 VGND VGND VPWR VPWR mem_addr[1] sky130_fd_sc_hd__buf_2
X_06017_ data_array.rdata0\[62\] net852 net1149 VGND VGND VPWR VPWR _03472_ sky130_fd_sc_hd__o21a_1
Xoutput252 net252 VGND VGND VPWR VPWR mem_addr[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput263 net263 VGND VGND VPWR VPWR mem_wdata[0] sky130_fd_sc_hd__buf_2
Xoutput274 net274 VGND VGND VPWR VPWR mem_wdata[1] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput285 net285 VGND VGND VPWR VPWR mem_wdata[2] sky130_fd_sc_hd__buf_2
XFILLER_0_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput296 net296 VGND VGND VPWR VPWR mem_wdata[3] sky130_fd_sc_hd__buf_2
XFILLER_181_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_250_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_250_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_114_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07968_ _05160_ _05161_ VGND VGND VPWR VPWR _00105_ sky130_fd_sc_hd__or2_1
XFILLER_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06919_ data_array.data0\[1\]\[16\] net1549 net1453 data_array.data0\[2\]\[16\] VGND
+ VGND VPWR VPWR _04208_ sky130_fd_sc_hd__a22o_1
X_09707_ net758 net3253 net611 VGND VGND VPWR VPWR _01459_ sky130_fd_sc_hd__mux2_1
X_07899_ data_array.data1\[0\]\[41\] net1335 net1241 data_array.data1\[3\]\[41\] _05098_
+ VGND VGND VPWR VPWR _05099_ sky130_fd_sc_hd__a221o_1
XFILLER_55_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_717 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09638_ net736 net3413 net615 VGND VGND VPWR VPWR _01390_ sky130_fd_sc_hd__mux2_1
XFILLER_130_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09569_ net1073 net2208 net399 VGND VGND VPWR VPWR _01321_ sky130_fd_sc_hd__mux2_1
X_11600_ clknet_leaf_140_clk _00408_ VGND VGND VPWR VPWR tag_array.tag1\[4\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12580_ clknet_leaf_154_clk _01274_ VGND VGND VPWR VPWR tag_array.tag0\[10\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_142_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11531_ clknet_leaf_175_clk _00339_ VGND VGND VPWR VPWR tag_array.valid1\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_12_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14250_ clknet_leaf_7_clk _02879_ VGND VGND VPWR VPWR data_array.data1\[12\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
X_11462_ clknet_leaf_2_clk _00272_ VGND VGND VPWR VPWR data_array.data0\[0\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13201_ clknet_leaf_77_clk _00095_ VGND VGND VPWR VPWR data_array.rdata1\[38\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_150_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10413_ net2251 net1000 net662 VGND VGND VPWR VPWR _02159_ sky130_fd_sc_hd__mux2_1
X_14181_ clknet_leaf_52_clk _02810_ VGND VGND VPWR VPWR data_array.data0\[2\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_11393_ clknet_leaf_132_clk _00203_ VGND VGND VPWR VPWR tag_array.tag1\[7\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_124_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_111_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13132_ clknet_leaf_106_clk _01826_ VGND VGND VPWR VPWR tag_array.tag0\[3\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_111_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10344_ net722 net3287 net592 VGND VGND VPWR VPWR _02091_ sky130_fd_sc_hd__mux2_1
XFILLER_98_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13063_ clknet_leaf_42_clk _01757_ VGND VGND VPWR VPWR data_array.data1\[13\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_140_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10275_ net2010 net1062 net641 VGND VGND VPWR VPWR _02022_ sky130_fd_sc_hd__mux2_1
XFILLER_151_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1400 _03513_ VGND VGND VPWR VPWR net1400 sky130_fd_sc_hd__buf_4
X_12014_ clknet_leaf_92_clk _00822_ VGND VGND VPWR VPWR data_array.data0\[6\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout1411 net1413 VGND VGND VPWR VPWR net1411 sky130_fd_sc_hd__clkbuf_4
Xfanout1422 _03513_ VGND VGND VPWR VPWR net1422 sky130_fd_sc_hd__clkbuf_4
Xfanout1433 net1434 VGND VGND VPWR VPWR net1433 sky130_fd_sc_hd__clkbuf_2
XFILLER_78_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_241_clk clknet_5_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_241_clk
+ sky130_fd_sc_hd__clkbuf_8
Xfanout1444 net1446 VGND VGND VPWR VPWR net1444 sky130_fd_sc_hd__clkbuf_4
Xfanout1455 net1458 VGND VGND VPWR VPWR net1455 sky130_fd_sc_hd__clkbuf_4
XFILLER_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1466 net1467 VGND VGND VPWR VPWR net1466 sky130_fd_sc_hd__clkbuf_4
Xfanout1477 net1495 VGND VGND VPWR VPWR net1477 sky130_fd_sc_hd__clkbuf_2
Xfanout490 net495 VGND VGND VPWR VPWR net490 sky130_fd_sc_hd__buf_4
Xfanout1488 net1495 VGND VGND VPWR VPWR net1488 sky130_fd_sc_hd__clkbuf_4
XFILLER_93_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1499 net1500 VGND VGND VPWR VPWR net1499 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13965_ clknet_leaf_198_clk _02594_ VGND VGND VPWR VPWR data_array.data1\[5\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12916_ clknet_leaf_127_clk _01610_ VGND VGND VPWR VPWR data_array.data0\[13\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_94_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13896_ clknet_leaf_227_clk _02525_ VGND VGND VPWR VPWR data_array.data1\[4\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_17_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12847_ clknet_leaf_63_clk _01541_ VGND VGND VPWR VPWR data_array.data0\[12\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_174_3711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12778_ clknet_leaf_158_clk _01472_ VGND VGND VPWR VPWR tag_array.tag0\[6\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_170_3619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11729_ clknet_leaf_169_clk _00537_ VGND VGND VPWR VPWR tag_array.tag0\[9\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14448_ clknet_leaf_265_clk _03071_ VGND VGND VPWR VPWR data_array.data1\[7\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_162_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold905 data_array.data0\[9\]\[11\] VGND VGND VPWR VPWR net2556 sky130_fd_sc_hd__dlygate4sd3_1
X_14379_ clknet_leaf_39_clk _03002_ VGND VGND VPWR VPWR data_array.data1\[10\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold916 data_array.data1\[13\]\[49\] VGND VGND VPWR VPWR net2567 sky130_fd_sc_hd__dlygate4sd3_1
Xhold927 tag_array.tag0\[14\]\[14\] VGND VGND VPWR VPWR net2578 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold938 data_array.data0\[14\]\[9\] VGND VGND VPWR VPWR net2589 sky130_fd_sc_hd__dlygate4sd3_1
Xhold949 tag_array.tag0\[6\]\[21\] VGND VGND VPWR VPWR net2600 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_142_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08940_ net1006 net2551 net428 VGND VGND VPWR VPWR _00696_ sky130_fd_sc_hd__mux2_1
XFILLER_131_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2306 tag_array.dirty0\[14\] VGND VGND VPWR VPWR net3957 sky130_fd_sc_hd__dlygate4sd3_1
X_08871_ net1020 net4531 net435 VGND VGND VPWR VPWR _00628_ sky130_fd_sc_hd__mux2_1
Xhold2317 data_array.data0\[15\]\[31\] VGND VGND VPWR VPWR net3968 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2328 data_array.data1\[12\]\[6\] VGND VGND VPWR VPWR net3979 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2339 tag_array.dirty0\[7\] VGND VGND VPWR VPWR net3990 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1605 lru_array.lru_mem\[10\] VGND VGND VPWR VPWR net3256 sky130_fd_sc_hd__dlygate4sd3_1
X_07822_ data_array.data1\[0\]\[34\] net1340 net1246 data_array.data1\[3\]\[34\] _05028_
+ VGND VGND VPWR VPWR _05029_ sky130_fd_sc_hd__a221o_1
XFILLER_57_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_232_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_232_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_9_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1616 tag_array.tag1\[14\]\[10\] VGND VGND VPWR VPWR net3267 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1627 data_array.data1\[5\]\[0\] VGND VGND VPWR VPWR net3278 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1638 tag_array.tag0\[12\]\[22\] VGND VGND VPWR VPWR net3289 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1649 data_array.data1\[9\]\[30\] VGND VGND VPWR VPWR net3300 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07753_ data_array.data1\[13\]\[28\] net1542 net1446 data_array.data1\[14\]\[28\]
+ VGND VGND VPWR VPWR _04966_ sky130_fd_sc_hd__a22o_1
X_06704_ tag_array.tag1\[13\]\[22\] net1552 net1456 tag_array.tag1\[14\]\[22\] VGND
+ VGND VPWR VPWR _04012_ sky130_fd_sc_hd__a22o_1
XFILLER_38_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07684_ data_array.data1\[8\]\[22\] net1348 net1254 data_array.data1\[11\]\[22\]
+ _04902_ VGND VGND VPWR VPWR _04903_ sky130_fd_sc_hd__a221o_1
XFILLER_25_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09423_ net975 net2423 net578 VGND VGND VPWR VPWR _01176_ sky130_fd_sc_hd__mux2_1
XFILLER_80_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06635_ net1633 _03943_ _03947_ net1207 VGND VGND VPWR VPWR _03950_ sky130_fd_sc_hd__a22o_1
XFILLER_80_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09354_ net987 net2485 net406 VGND VGND VPWR VPWR _01107_ sky130_fd_sc_hd__mux2_1
X_06566_ tag_array.tag1\[12\]\[9\] net1418 net1324 tag_array.tag1\[15\]\[9\] _03886_
+ VGND VGND VPWR VPWR _03887_ sky130_fd_sc_hd__a221o_1
XFILLER_80_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08305_ net1129 _05439_ VGND VGND VPWR VPWR _05440_ sky130_fd_sc_hd__and2_1
X_09285_ net741 net3558 net565 VGND VGND VPWR VPWR _01039_ sky130_fd_sc_hd__mux2_1
XFILLER_127_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06497_ tag_array.tag1\[5\]\[3\] net1561 net1465 tag_array.tag1\[6\]\[3\] VGND VGND
+ VPWR VPWR _03824_ sky130_fd_sc_hd__a22o_1
XFILLER_138_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08236_ _03140_ _03147_ VGND VGND VPWR VPWR _05392_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_95_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_706 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08167_ lru_array.lru_mem\[13\] net1564 net1468 lru_array.lru_mem\[14\] VGND VGND
+ VPWR VPWR _05342_ sky130_fd_sc_hd__a22o_1
XFILLER_134_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07118_ data_array.data0\[0\]\[34\] net1340 net1246 data_array.data0\[3\]\[34\] _04388_
+ VGND VGND VPWR VPWR _04389_ sky130_fd_sc_hd__a221o_1
XFILLER_118_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08098_ net1629 _05273_ _05277_ net1202 VGND VGND VPWR VPWR _05280_ sky130_fd_sc_hd__a22o_1
X_07049_ data_array.data0\[13\]\[28\] net1575 net1479 data_array.data0\[14\]\[28\]
+ VGND VGND VPWR VPWR _04326_ sky130_fd_sc_hd__a22o_1
XFILLER_0_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10060_ net784 net3655 net599 VGND VGND VPWR VPWR _01809_ sky130_fd_sc_hd__mux2_1
XFILLER_121_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_223_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_223_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_125_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2840 data_array.data1\[14\]\[1\] VGND VGND VPWR VPWR net4491 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2851 data_array.data0\[13\]\[27\] VGND VGND VPWR VPWR net4502 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2862 data_array.data1\[15\]\[42\] VGND VGND VPWR VPWR net4513 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2873 tag_array.tag0\[5\]\[8\] VGND VGND VPWR VPWR net4524 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_134_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2884 tag_array.tag1\[9\]\[15\] VGND VGND VPWR VPWR net4535 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2895 data_array.data0\[15\]\[46\] VGND VGND VPWR VPWR net4546 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_63_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10962_ net892 net4553 net528 VGND VGND VPWR VPWR _02707_ sky130_fd_sc_hd__mux2_1
X_13750_ clknet_leaf_261_clk _02379_ VGND VGND VPWR VPWR data_array.data1\[1\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
X_12701_ clknet_leaf_160_clk _01395_ VGND VGND VPWR VPWR tag_array.tag0\[8\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_43_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13681_ clknet_leaf_258_clk _02310_ VGND VGND VPWR VPWR data_array.data1\[15\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_67_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10893_ net915 net2861 net520 VGND VGND VPWR VPWR _02638_ sky130_fd_sc_hd__mux2_1
X_12632_ clknet_leaf_51_clk _01326_ VGND VGND VPWR VPWR data_array.data0\[15\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_84_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12563_ clknet_leaf_170_clk _01257_ VGND VGND VPWR VPWR tag_array.tag0\[11\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_180_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11514_ clknet_leaf_134_clk _00322_ VGND VGND VPWR VPWR tag_array.tag1\[9\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_14302_ clknet_leaf_24_clk _02931_ VGND VGND VPWR VPWR data_array.data1\[11\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_129_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12494_ clknet_leaf_244_clk _01188_ VGND VGND VPWR VPWR data_array.data1\[9\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14233_ clknet_leaf_250_clk _02862_ VGND VGND VPWR VPWR data_array.data1\[12\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_11445_ clknet_leaf_11_clk _00255_ VGND VGND VPWR VPWR data_array.data0\[0\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14164_ clknet_leaf_94_clk _02793_ VGND VGND VPWR VPWR data_array.data0\[2\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_11376_ net1647 net3957 net646 VGND VGND VPWR VPWR _03119_ sky130_fd_sc_hd__mux2_1
XFILLER_166_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_156_Right_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13115_ clknet_leaf_168_clk _01809_ VGND VGND VPWR VPWR tag_array.tag0\[3\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_10327_ net793 net3277 net592 VGND VGND VPWR VPWR _02074_ sky130_fd_sc_hd__mux2_1
XFILLER_125_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14095_ clknet_leaf_113_clk _02724_ VGND VGND VPWR VPWR data_array.data0\[1\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_79_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_167_3570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ clknet_leaf_206_clk _01740_ VGND VGND VPWR VPWR data_array.data0\[3\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
X_10258_ net712 net3377 net595 VGND VGND VPWR VPWR _02005_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_214_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_214_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_94_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1230 net1234 VGND VGND VPWR VPWR net1230 sky130_fd_sc_hd__buf_4
Xfanout1241 net1242 VGND VGND VPWR VPWR net1241 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_128_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10189_ net1049 net2295 net359 VGND VGND VPWR VPWR _01936_ sky130_fd_sc_hd__mux2_1
Xfanout1252 net1254 VGND VGND VPWR VPWR net1252 sky130_fd_sc_hd__clkbuf_4
XFILLER_121_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1263 net1264 VGND VGND VPWR VPWR net1263 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_163_3489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1274 net1276 VGND VGND VPWR VPWR net1274 sky130_fd_sc_hd__clkbuf_4
XFILLER_93_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1285 net1288 VGND VGND VPWR VPWR net1285 sky130_fd_sc_hd__clkbuf_4
Xfanout1296 net1298 VGND VGND VPWR VPWR net1296 sky130_fd_sc_hd__clkbuf_2
XFILLER_82_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13948_ clknet_leaf_211_clk _02577_ VGND VGND VPWR VPWR data_array.data1\[4\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_93_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13879_ clknet_leaf_78_clk _02508_ VGND VGND VPWR VPWR data_array.data1\[3\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06420_ tag_array.tag0\[5\]\[21\] net1598 net1502 tag_array.tag0\[6\]\[21\] VGND
+ VGND VPWR VPWR _03754_ sky130_fd_sc_hd__a22o_1
X_06351_ _03690_ _03691_ VGND VGND VPWR VPWR _00136_ sky130_fd_sc_hd__or2_1
XFILLER_30_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09070_ net1006 net2204 net412 VGND VGND VPWR VPWR _00824_ sky130_fd_sc_hd__mux2_1
X_06282_ tag_array.tag0\[4\]\[8\] net1409 net1315 tag_array.tag0\[7\]\[8\] _03628_
+ VGND VGND VPWR VPWR _03629_ sky130_fd_sc_hd__a221o_1
X_08021_ net1195 _05203_ _05207_ net1621 VGND VGND VPWR VPWR _05210_ sky130_fd_sc_hd__a22o_1
XFILLER_175_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold702 data_array.data0\[2\]\[55\] VGND VGND VPWR VPWR net2353 sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 data_array.data0\[9\]\[35\] VGND VGND VPWR VPWR net2364 sky130_fd_sc_hd__dlygate4sd3_1
Xhold724 tag_array.tag0\[10\]\[1\] VGND VGND VPWR VPWR net2375 sky130_fd_sc_hd__dlygate4sd3_1
Xhold735 data_array.data0\[14\]\[5\] VGND VGND VPWR VPWR net2386 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold746 tag_array.tag0\[2\]\[12\] VGND VGND VPWR VPWR net2397 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_157_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold757 tag_array.tag0\[10\]\[15\] VGND VGND VPWR VPWR net2408 sky130_fd_sc_hd__dlygate4sd3_1
Xhold768 data_array.data1\[0\]\[5\] VGND VGND VPWR VPWR net2419 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_123_Right_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold779 tag_array.tag0\[2\]\[0\] VGND VGND VPWR VPWR net2430 sky130_fd_sc_hd__dlygate4sd3_1
X_09972_ net941 net2542 net377 VGND VGND VPWR VPWR _01721_ sky130_fd_sc_hd__mux2_1
XFILLER_143_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08923_ net1072 net2471 net430 VGND VGND VPWR VPWR _00679_ sky130_fd_sc_hd__mux2_1
Xhold2103 data_array.data1\[9\]\[16\] VGND VGND VPWR VPWR net3754 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2114 tag_array.dirty0\[12\] VGND VGND VPWR VPWR net3765 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2125 data_array.data0\[7\]\[49\] VGND VGND VPWR VPWR net3776 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_205_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_205_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold2136 data_array.data0\[3\]\[28\] VGND VGND VPWR VPWR net3787 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1402 data_array.data0\[0\]\[0\] VGND VGND VPWR VPWR net3053 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2147 tag_array.tag0\[5\]\[13\] VGND VGND VPWR VPWR net3798 sky130_fd_sc_hd__dlygate4sd3_1
X_08854_ net1088 net3607 net436 VGND VGND VPWR VPWR _00611_ sky130_fd_sc_hd__mux2_1
Xhold2158 data_array.data0\[10\]\[51\] VGND VGND VPWR VPWR net3809 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1413 data_array.data0\[5\]\[4\] VGND VGND VPWR VPWR net3064 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1424 data_array.data1\[15\]\[30\] VGND VGND VPWR VPWR net3075 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2169 data_array.data1\[7\]\[57\] VGND VGND VPWR VPWR net3820 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1435 data_array.data1\[12\]\[33\] VGND VGND VPWR VPWR net3086 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07805_ data_array.data1\[12\]\[33\] net1398 net1304 data_array.data1\[15\]\[33\]
+ _05012_ VGND VGND VPWR VPWR _05013_ sky130_fd_sc_hd__a221o_1
Xhold1446 tag_array.tag0\[12\]\[24\] VGND VGND VPWR VPWR net3097 sky130_fd_sc_hd__dlygate4sd3_1
X_08785_ net3227 net1105 net442 VGND VGND VPWR VPWR _00543_ sky130_fd_sc_hd__mux2_1
XFILLER_57_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1457 data_array.data0\[15\]\[12\] VGND VGND VPWR VPWR net3108 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1468 data_array.data1\[3\]\[45\] VGND VGND VPWR VPWR net3119 sky130_fd_sc_hd__dlygate4sd3_1
X_05997_ data_array.rdata1\[55\] net835 net844 VGND VGND VPWR VPWR _03459_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_88_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1479 tag_array.tag1\[13\]\[22\] VGND VGND VPWR VPWR net3130 sky130_fd_sc_hd__dlygate4sd3_1
X_07736_ net1166 _04945_ _04949_ net1214 VGND VGND VPWR VPWR _04951_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_49_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07667_ data_array.data1\[1\]\[20\] net1605 net1509 data_array.data1\[2\]\[20\] VGND
+ VGND VPWR VPWR _04888_ sky130_fd_sc_hd__a22o_1
XFILLER_111_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09406_ net1041 net2309 net579 VGND VGND VPWR VPWR _01159_ sky130_fd_sc_hd__mux2_1
XFILLER_80_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06618_ tag_array.tag1\[1\]\[14\] net1558 net1462 tag_array.tag1\[2\]\[14\] VGND
+ VGND VPWR VPWR _03934_ sky130_fd_sc_hd__a22o_1
XFILLER_53_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07598_ data_array.data1\[4\]\[14\] net1379 net1285 data_array.data1\[7\]\[14\] _04824_
+ VGND VGND VPWR VPWR _04825_ sky130_fd_sc_hd__a221o_1
XFILLER_125_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06549_ _03870_ _03871_ VGND VGND VPWR VPWR _00178_ sky130_fd_sc_hd__or2_1
X_09337_ net1053 net4365 net406 VGND VGND VPWR VPWR _01090_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09268_ net706 net3319 net575 VGND VGND VPWR VPWR _01022_ sky130_fd_sc_hd__mux2_1
XFILLER_139_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08219_ fsm.tag_out1\[8\] net817 net809 fsm.tag_out0\[8\] _05380_ VGND VGND VPWR
+ VPWR _05381_ sky130_fd_sc_hd__a221o_1
XFILLER_14_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09199_ net785 net2355 net630 VGND VGND VPWR VPWR _00953_ sky130_fd_sc_hd__mux2_1
XFILLER_147_791 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11230_ net1110 net4503 net679 VGND VGND VPWR VPWR _02973_ sky130_fd_sc_hd__mux2_1
XFILLER_134_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11161_ net874 net4349 net548 VGND VGND VPWR VPWR _02904_ sky130_fd_sc_hd__mux2_1
XFILLER_20_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10112_ net1097 net4558 net366 VGND VGND VPWR VPWR _01860_ sky130_fd_sc_hd__mux2_1
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11092_ net2371 net895 net330 VGND VGND VPWR VPWR _02835_ sky130_fd_sc_hd__mux2_1
XFILLER_1_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10043_ net914 net2567 net561 VGND VGND VPWR VPWR _01792_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_145_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_959 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold51 tag_array.valid1\[14\] VGND VGND VPWR VPWR net1702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2670 data_array.data0\[5\]\[61\] VGND VGND VPWR VPWR net4321 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 tag_array.valid1\[4\] VGND VGND VPWR VPWR net1713 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_69_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2681 data_array.data1\[10\]\[2\] VGND VGND VPWR VPWR net4332 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 tag_array.valid1\[8\] VGND VGND VPWR VPWR net1724 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2692 data_array.data0\[3\]\[12\] VGND VGND VPWR VPWR net4343 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 data_array.data1\[0\]\[15\] VGND VGND VPWR VPWR net1735 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 data_array.data1\[2\]\[10\] VGND VGND VPWR VPWR net1746 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13802_ clknet_leaf_10_clk _02431_ VGND VGND VPWR VPWR data_array.data1\[2\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1980 data_array.data0\[15\]\[21\] VGND VGND VPWR VPWR net3631 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1991 tag_array.tag0\[1\]\[23\] VGND VGND VPWR VPWR net3642 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_21_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11994_ clknet_leaf_72_clk _00802_ VGND VGND VPWR VPWR data_array.data0\[6\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_962 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13733_ clknet_leaf_41_clk _02362_ VGND VGND VPWR VPWR data_array.data1\[1\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_10945_ net960 net2832 net528 VGND VGND VPWR VPWR _02690_ sky130_fd_sc_hd__mux2_1
XFILLER_16_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13664_ clknet_leaf_87_clk _02293_ VGND VGND VPWR VPWR data_array.data1\[15\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_10876_ net980 net4576 net514 VGND VGND VPWR VPWR _02621_ sky130_fd_sc_hd__mux2_1
X_12615_ clknet_leaf_190_clk _01309_ VGND VGND VPWR VPWR tag_array.tag0\[0\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_13595_ clknet_leaf_125_clk _02224_ VGND VGND VPWR VPWR data_array.data0\[9\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_157_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12546_ clknet_leaf_171_clk _01240_ VGND VGND VPWR VPWR tag_array.tag0\[11\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_77_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12477_ clknet_leaf_39_clk _01171_ VGND VGND VPWR VPWR data_array.data1\[9\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_169_3610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_4 _00101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14216_ clknet_leaf_174_clk _02845_ VGND VGND VPWR VPWR data_array.data1\[12\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_11428_ clknet_leaf_250_clk _00238_ VGND VGND VPWR VPWR data_array.data0\[0\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11359_ net858 net2236 net798 VGND VGND VPWR VPWR _03102_ sky130_fd_sc_hd__mux2_1
X_14147_ clknet_leaf_52_clk _02776_ VGND VGND VPWR VPWR data_array.data0\[1\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_165_3529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14078_ clknet_leaf_252_clk _02707_ VGND VGND VPWR VPWR data_array.data1\[6\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_140_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_5_Left_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_182_3854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05920_ net120 net1156 _03406_ _03407_ VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_182_3865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13029_ clknet_leaf_87_clk _01723_ VGND VGND VPWR VPWR data_array.data0\[3\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1060 net1061 VGND VGND VPWR VPWR net1060 sky130_fd_sc_hd__clkbuf_2
Xfanout1071 _05440_ VGND VGND VPWR VPWR net1071 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05851_ net159 net1150 _03360_ _03361_ VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__a22o_1
Xfanout1082 net1083 VGND VGND VPWR VPWR net1082 sky130_fd_sc_hd__clkbuf_2
Xfanout1093 _05428_ VGND VGND VPWR VPWR net1093 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08570_ net811 _05580_ VGND VGND VPWR VPWR _05600_ sky130_fd_sc_hd__and2_1
XFILLER_81_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05782_ net5 _03138_ _03271_ _03272_ _03298_ VGND VGND VPWR VPWR _03299_ sky130_fd_sc_hd__a2111o_1
XFILLER_148_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07521_ data_array.data1\[0\]\[7\] net1399 net1305 data_array.data1\[3\]\[7\] _04754_
+ VGND VGND VPWR VPWR _04755_ sky130_fd_sc_hd__a221o_1
XFILLER_179_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07452_ data_array.data1\[13\]\[1\] net1521 net1425 data_array.data1\[14\]\[1\] VGND
+ VGND VPWR VPWR _04692_ sky130_fd_sc_hd__a22o_1
XFILLER_34_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06403_ tag_array.tag0\[4\]\[19\] net1405 net1311 tag_array.tag0\[7\]\[19\] _03738_
+ VGND VGND VPWR VPWR _03739_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_44_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07383_ net1621 _04623_ _04627_ net1195 VGND VGND VPWR VPWR _04630_ sky130_fd_sc_hd__a22o_1
XFILLER_22_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09122_ net1054 net2784 net573 VGND VGND VPWR VPWR _00876_ sky130_fd_sc_hd__mux2_1
X_06334_ tag_array.tag0\[13\]\[13\] net1599 net1503 tag_array.tag0\[14\]\[13\] VGND
+ VGND VPWR VPWR _03676_ sky130_fd_sc_hd__a22o_1
XFILLER_124_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09053_ net1072 net2076 net414 VGND VGND VPWR VPWR _00807_ sky130_fd_sc_hd__mux2_1
XFILLER_175_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06265_ tag_array.tag0\[8\]\[7\] net1409 net1315 tag_array.tag0\[11\]\[7\] _03612_
+ VGND VGND VPWR VPWR _03613_ sky130_fd_sc_hd__a221o_1
XFILLER_163_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08004_ data_array.data1\[5\]\[51\] net1524 net1428 data_array.data1\[6\]\[51\] VGND
+ VGND VPWR VPWR _05194_ sky130_fd_sc_hd__a22o_1
Xhold510 data_array.data1\[4\]\[36\] VGND VGND VPWR VPWR net2161 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06196_ net1181 _03545_ _03549_ net1229 VGND VGND VPWR VPWR _03551_ sky130_fd_sc_hd__a22o_1
Xhold521 tag_array.tag1\[8\]\[1\] VGND VGND VPWR VPWR net2172 sky130_fd_sc_hd__dlygate4sd3_1
Xhold532 data_array.data1\[8\]\[15\] VGND VGND VPWR VPWR net2183 sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 tag_array.tag0\[15\]\[9\] VGND VGND VPWR VPWR net2194 sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 data_array.data0\[0\]\[55\] VGND VGND VPWR VPWR net2205 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold565 data_array.data1\[7\]\[2\] VGND VGND VPWR VPWR net2216 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_591 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold576 data_array.data1\[2\]\[0\] VGND VGND VPWR VPWR net2227 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold587 data_array.data1\[2\]\[44\] VGND VGND VPWR VPWR net2238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold598 tag_array.tag0\[15\]\[20\] VGND VGND VPWR VPWR net2249 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09955_ net1010 net3007 net370 VGND VGND VPWR VPWR _01704_ sky130_fd_sc_hd__mux2_1
XFILLER_106_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_5_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08906_ net881 net4591 net437 VGND VGND VPWR VPWR _00663_ sky130_fd_sc_hd__mux2_1
X_09886_ net926 net4407 net378 VGND VGND VPWR VPWR _01636_ sky130_fd_sc_hd__mux2_1
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1210 data_array.data1\[5\]\[49\] VGND VGND VPWR VPWR net2861 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1221 data_array.data0\[11\]\[36\] VGND VGND VPWR VPWR net2872 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1232 data_array.data0\[3\]\[8\] VGND VGND VPWR VPWR net2883 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08837_ net2475 net897 net442 VGND VGND VPWR VPWR _00595_ sky130_fd_sc_hd__mux2_1
Xhold1243 data_array.data1\[5\]\[22\] VGND VGND VPWR VPWR net2894 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1254 tag_array.tag0\[2\]\[23\] VGND VGND VPWR VPWR net2905 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1265 data_array.data0\[8\]\[26\] VGND VGND VPWR VPWR net2916 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1276 data_array.data1\[13\]\[19\] VGND VGND VPWR VPWR net2927 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1287 data_array.data1\[10\]\[56\] VGND VGND VPWR VPWR net2938 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1298 tag_array.tag1\[12\]\[7\] VGND VGND VPWR VPWR net2949 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08768_ net752 net2692 net451 VGND VGND VPWR VPWR _00527_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_140_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07719_ data_array.data1\[0\]\[25\] net1329 net1235 data_array.data1\[3\]\[25\] _04934_
+ VGND VGND VPWR VPWR _04935_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_64_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08699_ net1733 net728 net487 VGND VGND VPWR VPWR _00458_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10730_ net1054 net4451 net496 VGND VGND VPWR VPWR _02475_ sky130_fd_sc_hd__mux2_1
XFILLER_14_848 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10661_ net2206 net1074 net484 VGND VGND VPWR VPWR _02406_ sky130_fd_sc_hd__mux2_1
XFILLER_139_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12400_ clknet_leaf_15_clk _01094_ VGND VGND VPWR VPWR data_array.data0\[14\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_13380_ clknet_leaf_174_clk _02010_ VGND VGND VPWR VPWR data_array.data1\[8\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_10592_ net1903 net1094 net472 VGND VGND VPWR VPWR _02337_ sky130_fd_sc_hd__mux2_1
XFILLER_167_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12331_ clknet_leaf_201_clk _00004_ VGND VGND VPWR VPWR data_array.rdata0\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_126_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12262_ clknet_leaf_95_clk _01020_ VGND VGND VPWR VPWR tag_array.tag1\[14\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_79_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_366 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11213_ net922 net4391 net657 VGND VGND VPWR VPWR _02956_ sky130_fd_sc_hd__mux2_1
X_14001_ clknet_leaf_258_clk _02630_ VGND VGND VPWR VPWR data_array.data1\[5\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_107_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12193_ clknet_leaf_145_clk _00131_ VGND VGND VPWR VPWR fsm.tag_out0\[0\] sky130_fd_sc_hd__dfxtp_2
X_11144_ net943 net3073 net550 VGND VGND VPWR VPWR _02887_ sky130_fd_sc_hd__mux2_1
XFILLER_1_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11075_ net1889 net961 net330 VGND VGND VPWR VPWR _02818_ sky130_fd_sc_hd__mux2_1
XFILLER_1_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput130 mem_rdata[38] VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_1
Xinput141 mem_rdata[48] VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10026_ net980 net3132 net554 VGND VGND VPWR VPWR _01775_ sky130_fd_sc_hd__mux2_1
Xinput152 mem_rdata[58] VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_160_3437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput163 mem_ready VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_2
XFILLER_63_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11977_ clknet_leaf_1_clk _00785_ VGND VGND VPWR VPWR data_array.data0\[4\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13716_ clknet_leaf_85_clk _02345_ VGND VGND VPWR VPWR data_array.data1\[1\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_10928_ net1030 net3310 net536 VGND VGND VPWR VPWR _02673_ sky130_fd_sc_hd__mux2_1
XFILLER_60_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13647_ clknet_leaf_82_clk _02276_ VGND VGND VPWR VPWR data_array.data1\[15\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_158_3399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10859_ net1049 net1955 net520 VGND VGND VPWR VPWR _02604_ sky130_fd_sc_hd__mux2_1
XFILLER_31_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13578_ clknet_leaf_47_clk _02207_ VGND VGND VPWR VPWR data_array.data0\[9\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_145_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12529_ clknet_leaf_32_clk _01223_ VGND VGND VPWR VPWR tag_array.tag1\[11\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_157_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06050_ fsm.tag_out0\[7\] net1121 _03488_ VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_10_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_184_3905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_184_3916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09740_ net728 net2186 net683 VGND VGND VPWR VPWR _01492_ sky130_fd_sc_hd__mux2_1
X_06952_ data_array.data0\[1\]\[19\] net1582 net1486 data_array.data0\[2\]\[19\] VGND
+ VGND VPWR VPWR _04238_ sky130_fd_sc_hd__a22o_1
XFILLER_100_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
.ends

