module cache_controller (clk,
    cpu_read,
    cpu_ready,
    cpu_write,
    mem_read,
    mem_ready,
    mem_write,
    reset,
    cpu_addr,
    cpu_rdata,
    cpu_wdata,
    mem_addr,
    mem_rdata,
    mem_wdata);
 input clk;
 input cpu_read;
 output cpu_ready;
 input cpu_write;
 output mem_read;
 input mem_ready;
 output mem_write;
 input reset;
 input [31:0] cpu_addr;
 output [63:0] cpu_rdata;
 input [63:0] cpu_wdata;
 output [31:0] mem_addr;
 input [63:0] mem_rdata;
 output [63:0] mem_wdata;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire \data_array.data0[0][0] ;
 wire \data_array.data0[0][10] ;
 wire \data_array.data0[0][11] ;
 wire \data_array.data0[0][12] ;
 wire \data_array.data0[0][13] ;
 wire \data_array.data0[0][14] ;
 wire \data_array.data0[0][15] ;
 wire \data_array.data0[0][16] ;
 wire \data_array.data0[0][17] ;
 wire \data_array.data0[0][18] ;
 wire \data_array.data0[0][19] ;
 wire \data_array.data0[0][1] ;
 wire \data_array.data0[0][20] ;
 wire \data_array.data0[0][21] ;
 wire \data_array.data0[0][22] ;
 wire \data_array.data0[0][23] ;
 wire \data_array.data0[0][24] ;
 wire \data_array.data0[0][25] ;
 wire \data_array.data0[0][26] ;
 wire \data_array.data0[0][27] ;
 wire \data_array.data0[0][28] ;
 wire \data_array.data0[0][29] ;
 wire \data_array.data0[0][2] ;
 wire \data_array.data0[0][30] ;
 wire \data_array.data0[0][31] ;
 wire \data_array.data0[0][32] ;
 wire \data_array.data0[0][33] ;
 wire \data_array.data0[0][34] ;
 wire \data_array.data0[0][35] ;
 wire \data_array.data0[0][36] ;
 wire \data_array.data0[0][37] ;
 wire \data_array.data0[0][38] ;
 wire \data_array.data0[0][39] ;
 wire \data_array.data0[0][3] ;
 wire \data_array.data0[0][40] ;
 wire \data_array.data0[0][41] ;
 wire \data_array.data0[0][42] ;
 wire \data_array.data0[0][43] ;
 wire \data_array.data0[0][44] ;
 wire \data_array.data0[0][45] ;
 wire \data_array.data0[0][46] ;
 wire \data_array.data0[0][47] ;
 wire \data_array.data0[0][48] ;
 wire \data_array.data0[0][49] ;
 wire \data_array.data0[0][4] ;
 wire \data_array.data0[0][50] ;
 wire \data_array.data0[0][51] ;
 wire \data_array.data0[0][52] ;
 wire \data_array.data0[0][53] ;
 wire \data_array.data0[0][54] ;
 wire \data_array.data0[0][55] ;
 wire \data_array.data0[0][56] ;
 wire \data_array.data0[0][57] ;
 wire \data_array.data0[0][58] ;
 wire \data_array.data0[0][59] ;
 wire \data_array.data0[0][5] ;
 wire \data_array.data0[0][60] ;
 wire \data_array.data0[0][61] ;
 wire \data_array.data0[0][62] ;
 wire \data_array.data0[0][63] ;
 wire \data_array.data0[0][6] ;
 wire \data_array.data0[0][7] ;
 wire \data_array.data0[0][8] ;
 wire \data_array.data0[0][9] ;
 wire \data_array.data0[10][0] ;
 wire \data_array.data0[10][10] ;
 wire \data_array.data0[10][11] ;
 wire \data_array.data0[10][12] ;
 wire \data_array.data0[10][13] ;
 wire \data_array.data0[10][14] ;
 wire \data_array.data0[10][15] ;
 wire \data_array.data0[10][16] ;
 wire \data_array.data0[10][17] ;
 wire \data_array.data0[10][18] ;
 wire \data_array.data0[10][19] ;
 wire \data_array.data0[10][1] ;
 wire \data_array.data0[10][20] ;
 wire \data_array.data0[10][21] ;
 wire \data_array.data0[10][22] ;
 wire \data_array.data0[10][23] ;
 wire \data_array.data0[10][24] ;
 wire \data_array.data0[10][25] ;
 wire \data_array.data0[10][26] ;
 wire \data_array.data0[10][27] ;
 wire \data_array.data0[10][28] ;
 wire \data_array.data0[10][29] ;
 wire \data_array.data0[10][2] ;
 wire \data_array.data0[10][30] ;
 wire \data_array.data0[10][31] ;
 wire \data_array.data0[10][32] ;
 wire \data_array.data0[10][33] ;
 wire \data_array.data0[10][34] ;
 wire \data_array.data0[10][35] ;
 wire \data_array.data0[10][36] ;
 wire \data_array.data0[10][37] ;
 wire \data_array.data0[10][38] ;
 wire \data_array.data0[10][39] ;
 wire \data_array.data0[10][3] ;
 wire \data_array.data0[10][40] ;
 wire \data_array.data0[10][41] ;
 wire \data_array.data0[10][42] ;
 wire \data_array.data0[10][43] ;
 wire \data_array.data0[10][44] ;
 wire \data_array.data0[10][45] ;
 wire \data_array.data0[10][46] ;
 wire \data_array.data0[10][47] ;
 wire \data_array.data0[10][48] ;
 wire \data_array.data0[10][49] ;
 wire \data_array.data0[10][4] ;
 wire \data_array.data0[10][50] ;
 wire \data_array.data0[10][51] ;
 wire \data_array.data0[10][52] ;
 wire \data_array.data0[10][53] ;
 wire \data_array.data0[10][54] ;
 wire \data_array.data0[10][55] ;
 wire \data_array.data0[10][56] ;
 wire \data_array.data0[10][57] ;
 wire \data_array.data0[10][58] ;
 wire \data_array.data0[10][59] ;
 wire \data_array.data0[10][5] ;
 wire \data_array.data0[10][60] ;
 wire \data_array.data0[10][61] ;
 wire \data_array.data0[10][62] ;
 wire \data_array.data0[10][63] ;
 wire \data_array.data0[10][6] ;
 wire \data_array.data0[10][7] ;
 wire \data_array.data0[10][8] ;
 wire \data_array.data0[10][9] ;
 wire \data_array.data0[11][0] ;
 wire \data_array.data0[11][10] ;
 wire \data_array.data0[11][11] ;
 wire \data_array.data0[11][12] ;
 wire \data_array.data0[11][13] ;
 wire \data_array.data0[11][14] ;
 wire \data_array.data0[11][15] ;
 wire \data_array.data0[11][16] ;
 wire \data_array.data0[11][17] ;
 wire \data_array.data0[11][18] ;
 wire \data_array.data0[11][19] ;
 wire \data_array.data0[11][1] ;
 wire \data_array.data0[11][20] ;
 wire \data_array.data0[11][21] ;
 wire \data_array.data0[11][22] ;
 wire \data_array.data0[11][23] ;
 wire \data_array.data0[11][24] ;
 wire \data_array.data0[11][25] ;
 wire \data_array.data0[11][26] ;
 wire \data_array.data0[11][27] ;
 wire \data_array.data0[11][28] ;
 wire \data_array.data0[11][29] ;
 wire \data_array.data0[11][2] ;
 wire \data_array.data0[11][30] ;
 wire \data_array.data0[11][31] ;
 wire \data_array.data0[11][32] ;
 wire \data_array.data0[11][33] ;
 wire \data_array.data0[11][34] ;
 wire \data_array.data0[11][35] ;
 wire \data_array.data0[11][36] ;
 wire \data_array.data0[11][37] ;
 wire \data_array.data0[11][38] ;
 wire \data_array.data0[11][39] ;
 wire \data_array.data0[11][3] ;
 wire \data_array.data0[11][40] ;
 wire \data_array.data0[11][41] ;
 wire \data_array.data0[11][42] ;
 wire \data_array.data0[11][43] ;
 wire \data_array.data0[11][44] ;
 wire \data_array.data0[11][45] ;
 wire \data_array.data0[11][46] ;
 wire \data_array.data0[11][47] ;
 wire \data_array.data0[11][48] ;
 wire \data_array.data0[11][49] ;
 wire \data_array.data0[11][4] ;
 wire \data_array.data0[11][50] ;
 wire \data_array.data0[11][51] ;
 wire \data_array.data0[11][52] ;
 wire \data_array.data0[11][53] ;
 wire \data_array.data0[11][54] ;
 wire \data_array.data0[11][55] ;
 wire \data_array.data0[11][56] ;
 wire \data_array.data0[11][57] ;
 wire \data_array.data0[11][58] ;
 wire \data_array.data0[11][59] ;
 wire \data_array.data0[11][5] ;
 wire \data_array.data0[11][60] ;
 wire \data_array.data0[11][61] ;
 wire \data_array.data0[11][62] ;
 wire \data_array.data0[11][63] ;
 wire \data_array.data0[11][6] ;
 wire \data_array.data0[11][7] ;
 wire \data_array.data0[11][8] ;
 wire \data_array.data0[11][9] ;
 wire \data_array.data0[12][0] ;
 wire \data_array.data0[12][10] ;
 wire \data_array.data0[12][11] ;
 wire \data_array.data0[12][12] ;
 wire \data_array.data0[12][13] ;
 wire \data_array.data0[12][14] ;
 wire \data_array.data0[12][15] ;
 wire \data_array.data0[12][16] ;
 wire \data_array.data0[12][17] ;
 wire \data_array.data0[12][18] ;
 wire \data_array.data0[12][19] ;
 wire \data_array.data0[12][1] ;
 wire \data_array.data0[12][20] ;
 wire \data_array.data0[12][21] ;
 wire \data_array.data0[12][22] ;
 wire \data_array.data0[12][23] ;
 wire \data_array.data0[12][24] ;
 wire \data_array.data0[12][25] ;
 wire \data_array.data0[12][26] ;
 wire \data_array.data0[12][27] ;
 wire \data_array.data0[12][28] ;
 wire \data_array.data0[12][29] ;
 wire \data_array.data0[12][2] ;
 wire \data_array.data0[12][30] ;
 wire \data_array.data0[12][31] ;
 wire \data_array.data0[12][32] ;
 wire \data_array.data0[12][33] ;
 wire \data_array.data0[12][34] ;
 wire \data_array.data0[12][35] ;
 wire \data_array.data0[12][36] ;
 wire \data_array.data0[12][37] ;
 wire \data_array.data0[12][38] ;
 wire \data_array.data0[12][39] ;
 wire \data_array.data0[12][3] ;
 wire \data_array.data0[12][40] ;
 wire \data_array.data0[12][41] ;
 wire \data_array.data0[12][42] ;
 wire \data_array.data0[12][43] ;
 wire \data_array.data0[12][44] ;
 wire \data_array.data0[12][45] ;
 wire \data_array.data0[12][46] ;
 wire \data_array.data0[12][47] ;
 wire \data_array.data0[12][48] ;
 wire \data_array.data0[12][49] ;
 wire \data_array.data0[12][4] ;
 wire \data_array.data0[12][50] ;
 wire \data_array.data0[12][51] ;
 wire \data_array.data0[12][52] ;
 wire \data_array.data0[12][53] ;
 wire \data_array.data0[12][54] ;
 wire \data_array.data0[12][55] ;
 wire \data_array.data0[12][56] ;
 wire \data_array.data0[12][57] ;
 wire \data_array.data0[12][58] ;
 wire \data_array.data0[12][59] ;
 wire \data_array.data0[12][5] ;
 wire \data_array.data0[12][60] ;
 wire \data_array.data0[12][61] ;
 wire \data_array.data0[12][62] ;
 wire \data_array.data0[12][63] ;
 wire \data_array.data0[12][6] ;
 wire \data_array.data0[12][7] ;
 wire \data_array.data0[12][8] ;
 wire \data_array.data0[12][9] ;
 wire \data_array.data0[13][0] ;
 wire \data_array.data0[13][10] ;
 wire \data_array.data0[13][11] ;
 wire \data_array.data0[13][12] ;
 wire \data_array.data0[13][13] ;
 wire \data_array.data0[13][14] ;
 wire \data_array.data0[13][15] ;
 wire \data_array.data0[13][16] ;
 wire \data_array.data0[13][17] ;
 wire \data_array.data0[13][18] ;
 wire \data_array.data0[13][19] ;
 wire \data_array.data0[13][1] ;
 wire \data_array.data0[13][20] ;
 wire \data_array.data0[13][21] ;
 wire \data_array.data0[13][22] ;
 wire \data_array.data0[13][23] ;
 wire \data_array.data0[13][24] ;
 wire \data_array.data0[13][25] ;
 wire \data_array.data0[13][26] ;
 wire \data_array.data0[13][27] ;
 wire \data_array.data0[13][28] ;
 wire \data_array.data0[13][29] ;
 wire \data_array.data0[13][2] ;
 wire \data_array.data0[13][30] ;
 wire \data_array.data0[13][31] ;
 wire \data_array.data0[13][32] ;
 wire \data_array.data0[13][33] ;
 wire \data_array.data0[13][34] ;
 wire \data_array.data0[13][35] ;
 wire \data_array.data0[13][36] ;
 wire \data_array.data0[13][37] ;
 wire \data_array.data0[13][38] ;
 wire \data_array.data0[13][39] ;
 wire \data_array.data0[13][3] ;
 wire \data_array.data0[13][40] ;
 wire \data_array.data0[13][41] ;
 wire \data_array.data0[13][42] ;
 wire \data_array.data0[13][43] ;
 wire \data_array.data0[13][44] ;
 wire \data_array.data0[13][45] ;
 wire \data_array.data0[13][46] ;
 wire \data_array.data0[13][47] ;
 wire \data_array.data0[13][48] ;
 wire \data_array.data0[13][49] ;
 wire \data_array.data0[13][4] ;
 wire \data_array.data0[13][50] ;
 wire \data_array.data0[13][51] ;
 wire \data_array.data0[13][52] ;
 wire \data_array.data0[13][53] ;
 wire \data_array.data0[13][54] ;
 wire \data_array.data0[13][55] ;
 wire \data_array.data0[13][56] ;
 wire \data_array.data0[13][57] ;
 wire \data_array.data0[13][58] ;
 wire \data_array.data0[13][59] ;
 wire \data_array.data0[13][5] ;
 wire \data_array.data0[13][60] ;
 wire \data_array.data0[13][61] ;
 wire \data_array.data0[13][62] ;
 wire \data_array.data0[13][63] ;
 wire \data_array.data0[13][6] ;
 wire \data_array.data0[13][7] ;
 wire \data_array.data0[13][8] ;
 wire \data_array.data0[13][9] ;
 wire \data_array.data0[14][0] ;
 wire \data_array.data0[14][10] ;
 wire \data_array.data0[14][11] ;
 wire \data_array.data0[14][12] ;
 wire \data_array.data0[14][13] ;
 wire \data_array.data0[14][14] ;
 wire \data_array.data0[14][15] ;
 wire \data_array.data0[14][16] ;
 wire \data_array.data0[14][17] ;
 wire \data_array.data0[14][18] ;
 wire \data_array.data0[14][19] ;
 wire \data_array.data0[14][1] ;
 wire \data_array.data0[14][20] ;
 wire \data_array.data0[14][21] ;
 wire \data_array.data0[14][22] ;
 wire \data_array.data0[14][23] ;
 wire \data_array.data0[14][24] ;
 wire \data_array.data0[14][25] ;
 wire \data_array.data0[14][26] ;
 wire \data_array.data0[14][27] ;
 wire \data_array.data0[14][28] ;
 wire \data_array.data0[14][29] ;
 wire \data_array.data0[14][2] ;
 wire \data_array.data0[14][30] ;
 wire \data_array.data0[14][31] ;
 wire \data_array.data0[14][32] ;
 wire \data_array.data0[14][33] ;
 wire \data_array.data0[14][34] ;
 wire \data_array.data0[14][35] ;
 wire \data_array.data0[14][36] ;
 wire \data_array.data0[14][37] ;
 wire \data_array.data0[14][38] ;
 wire \data_array.data0[14][39] ;
 wire \data_array.data0[14][3] ;
 wire \data_array.data0[14][40] ;
 wire \data_array.data0[14][41] ;
 wire \data_array.data0[14][42] ;
 wire \data_array.data0[14][43] ;
 wire \data_array.data0[14][44] ;
 wire \data_array.data0[14][45] ;
 wire \data_array.data0[14][46] ;
 wire \data_array.data0[14][47] ;
 wire \data_array.data0[14][48] ;
 wire \data_array.data0[14][49] ;
 wire \data_array.data0[14][4] ;
 wire \data_array.data0[14][50] ;
 wire \data_array.data0[14][51] ;
 wire \data_array.data0[14][52] ;
 wire \data_array.data0[14][53] ;
 wire \data_array.data0[14][54] ;
 wire \data_array.data0[14][55] ;
 wire \data_array.data0[14][56] ;
 wire \data_array.data0[14][57] ;
 wire \data_array.data0[14][58] ;
 wire \data_array.data0[14][59] ;
 wire \data_array.data0[14][5] ;
 wire \data_array.data0[14][60] ;
 wire \data_array.data0[14][61] ;
 wire \data_array.data0[14][62] ;
 wire \data_array.data0[14][63] ;
 wire \data_array.data0[14][6] ;
 wire \data_array.data0[14][7] ;
 wire \data_array.data0[14][8] ;
 wire \data_array.data0[14][9] ;
 wire \data_array.data0[15][0] ;
 wire \data_array.data0[15][10] ;
 wire \data_array.data0[15][11] ;
 wire \data_array.data0[15][12] ;
 wire \data_array.data0[15][13] ;
 wire \data_array.data0[15][14] ;
 wire \data_array.data0[15][15] ;
 wire \data_array.data0[15][16] ;
 wire \data_array.data0[15][17] ;
 wire \data_array.data0[15][18] ;
 wire \data_array.data0[15][19] ;
 wire \data_array.data0[15][1] ;
 wire \data_array.data0[15][20] ;
 wire \data_array.data0[15][21] ;
 wire \data_array.data0[15][22] ;
 wire \data_array.data0[15][23] ;
 wire \data_array.data0[15][24] ;
 wire \data_array.data0[15][25] ;
 wire \data_array.data0[15][26] ;
 wire \data_array.data0[15][27] ;
 wire \data_array.data0[15][28] ;
 wire \data_array.data0[15][29] ;
 wire \data_array.data0[15][2] ;
 wire \data_array.data0[15][30] ;
 wire \data_array.data0[15][31] ;
 wire \data_array.data0[15][32] ;
 wire \data_array.data0[15][33] ;
 wire \data_array.data0[15][34] ;
 wire \data_array.data0[15][35] ;
 wire \data_array.data0[15][36] ;
 wire \data_array.data0[15][37] ;
 wire \data_array.data0[15][38] ;
 wire \data_array.data0[15][39] ;
 wire \data_array.data0[15][3] ;
 wire \data_array.data0[15][40] ;
 wire \data_array.data0[15][41] ;
 wire \data_array.data0[15][42] ;
 wire \data_array.data0[15][43] ;
 wire \data_array.data0[15][44] ;
 wire \data_array.data0[15][45] ;
 wire \data_array.data0[15][46] ;
 wire \data_array.data0[15][47] ;
 wire \data_array.data0[15][48] ;
 wire \data_array.data0[15][49] ;
 wire \data_array.data0[15][4] ;
 wire \data_array.data0[15][50] ;
 wire \data_array.data0[15][51] ;
 wire \data_array.data0[15][52] ;
 wire \data_array.data0[15][53] ;
 wire \data_array.data0[15][54] ;
 wire \data_array.data0[15][55] ;
 wire \data_array.data0[15][56] ;
 wire \data_array.data0[15][57] ;
 wire \data_array.data0[15][58] ;
 wire \data_array.data0[15][59] ;
 wire \data_array.data0[15][5] ;
 wire \data_array.data0[15][60] ;
 wire \data_array.data0[15][61] ;
 wire \data_array.data0[15][62] ;
 wire \data_array.data0[15][63] ;
 wire \data_array.data0[15][6] ;
 wire \data_array.data0[15][7] ;
 wire \data_array.data0[15][8] ;
 wire \data_array.data0[15][9] ;
 wire \data_array.data0[1][0] ;
 wire \data_array.data0[1][10] ;
 wire \data_array.data0[1][11] ;
 wire \data_array.data0[1][12] ;
 wire \data_array.data0[1][13] ;
 wire \data_array.data0[1][14] ;
 wire \data_array.data0[1][15] ;
 wire \data_array.data0[1][16] ;
 wire \data_array.data0[1][17] ;
 wire \data_array.data0[1][18] ;
 wire \data_array.data0[1][19] ;
 wire \data_array.data0[1][1] ;
 wire \data_array.data0[1][20] ;
 wire \data_array.data0[1][21] ;
 wire \data_array.data0[1][22] ;
 wire \data_array.data0[1][23] ;
 wire \data_array.data0[1][24] ;
 wire \data_array.data0[1][25] ;
 wire \data_array.data0[1][26] ;
 wire \data_array.data0[1][27] ;
 wire \data_array.data0[1][28] ;
 wire \data_array.data0[1][29] ;
 wire \data_array.data0[1][2] ;
 wire \data_array.data0[1][30] ;
 wire \data_array.data0[1][31] ;
 wire \data_array.data0[1][32] ;
 wire \data_array.data0[1][33] ;
 wire \data_array.data0[1][34] ;
 wire \data_array.data0[1][35] ;
 wire \data_array.data0[1][36] ;
 wire \data_array.data0[1][37] ;
 wire \data_array.data0[1][38] ;
 wire \data_array.data0[1][39] ;
 wire \data_array.data0[1][3] ;
 wire \data_array.data0[1][40] ;
 wire \data_array.data0[1][41] ;
 wire \data_array.data0[1][42] ;
 wire \data_array.data0[1][43] ;
 wire \data_array.data0[1][44] ;
 wire \data_array.data0[1][45] ;
 wire \data_array.data0[1][46] ;
 wire \data_array.data0[1][47] ;
 wire \data_array.data0[1][48] ;
 wire \data_array.data0[1][49] ;
 wire \data_array.data0[1][4] ;
 wire \data_array.data0[1][50] ;
 wire \data_array.data0[1][51] ;
 wire \data_array.data0[1][52] ;
 wire \data_array.data0[1][53] ;
 wire \data_array.data0[1][54] ;
 wire \data_array.data0[1][55] ;
 wire \data_array.data0[1][56] ;
 wire \data_array.data0[1][57] ;
 wire \data_array.data0[1][58] ;
 wire \data_array.data0[1][59] ;
 wire \data_array.data0[1][5] ;
 wire \data_array.data0[1][60] ;
 wire \data_array.data0[1][61] ;
 wire \data_array.data0[1][62] ;
 wire \data_array.data0[1][63] ;
 wire \data_array.data0[1][6] ;
 wire \data_array.data0[1][7] ;
 wire \data_array.data0[1][8] ;
 wire \data_array.data0[1][9] ;
 wire \data_array.data0[2][0] ;
 wire \data_array.data0[2][10] ;
 wire \data_array.data0[2][11] ;
 wire \data_array.data0[2][12] ;
 wire \data_array.data0[2][13] ;
 wire \data_array.data0[2][14] ;
 wire \data_array.data0[2][15] ;
 wire \data_array.data0[2][16] ;
 wire \data_array.data0[2][17] ;
 wire \data_array.data0[2][18] ;
 wire \data_array.data0[2][19] ;
 wire \data_array.data0[2][1] ;
 wire \data_array.data0[2][20] ;
 wire \data_array.data0[2][21] ;
 wire \data_array.data0[2][22] ;
 wire \data_array.data0[2][23] ;
 wire \data_array.data0[2][24] ;
 wire \data_array.data0[2][25] ;
 wire \data_array.data0[2][26] ;
 wire \data_array.data0[2][27] ;
 wire \data_array.data0[2][28] ;
 wire \data_array.data0[2][29] ;
 wire \data_array.data0[2][2] ;
 wire \data_array.data0[2][30] ;
 wire \data_array.data0[2][31] ;
 wire \data_array.data0[2][32] ;
 wire \data_array.data0[2][33] ;
 wire \data_array.data0[2][34] ;
 wire \data_array.data0[2][35] ;
 wire \data_array.data0[2][36] ;
 wire \data_array.data0[2][37] ;
 wire \data_array.data0[2][38] ;
 wire \data_array.data0[2][39] ;
 wire \data_array.data0[2][3] ;
 wire \data_array.data0[2][40] ;
 wire \data_array.data0[2][41] ;
 wire \data_array.data0[2][42] ;
 wire \data_array.data0[2][43] ;
 wire \data_array.data0[2][44] ;
 wire \data_array.data0[2][45] ;
 wire \data_array.data0[2][46] ;
 wire \data_array.data0[2][47] ;
 wire \data_array.data0[2][48] ;
 wire \data_array.data0[2][49] ;
 wire \data_array.data0[2][4] ;
 wire \data_array.data0[2][50] ;
 wire \data_array.data0[2][51] ;
 wire \data_array.data0[2][52] ;
 wire \data_array.data0[2][53] ;
 wire \data_array.data0[2][54] ;
 wire \data_array.data0[2][55] ;
 wire \data_array.data0[2][56] ;
 wire \data_array.data0[2][57] ;
 wire \data_array.data0[2][58] ;
 wire \data_array.data0[2][59] ;
 wire \data_array.data0[2][5] ;
 wire \data_array.data0[2][60] ;
 wire \data_array.data0[2][61] ;
 wire \data_array.data0[2][62] ;
 wire \data_array.data0[2][63] ;
 wire \data_array.data0[2][6] ;
 wire \data_array.data0[2][7] ;
 wire \data_array.data0[2][8] ;
 wire \data_array.data0[2][9] ;
 wire \data_array.data0[3][0] ;
 wire \data_array.data0[3][10] ;
 wire \data_array.data0[3][11] ;
 wire \data_array.data0[3][12] ;
 wire \data_array.data0[3][13] ;
 wire \data_array.data0[3][14] ;
 wire \data_array.data0[3][15] ;
 wire \data_array.data0[3][16] ;
 wire \data_array.data0[3][17] ;
 wire \data_array.data0[3][18] ;
 wire \data_array.data0[3][19] ;
 wire \data_array.data0[3][1] ;
 wire \data_array.data0[3][20] ;
 wire \data_array.data0[3][21] ;
 wire \data_array.data0[3][22] ;
 wire \data_array.data0[3][23] ;
 wire \data_array.data0[3][24] ;
 wire \data_array.data0[3][25] ;
 wire \data_array.data0[3][26] ;
 wire \data_array.data0[3][27] ;
 wire \data_array.data0[3][28] ;
 wire \data_array.data0[3][29] ;
 wire \data_array.data0[3][2] ;
 wire \data_array.data0[3][30] ;
 wire \data_array.data0[3][31] ;
 wire \data_array.data0[3][32] ;
 wire \data_array.data0[3][33] ;
 wire \data_array.data0[3][34] ;
 wire \data_array.data0[3][35] ;
 wire \data_array.data0[3][36] ;
 wire \data_array.data0[3][37] ;
 wire \data_array.data0[3][38] ;
 wire \data_array.data0[3][39] ;
 wire \data_array.data0[3][3] ;
 wire \data_array.data0[3][40] ;
 wire \data_array.data0[3][41] ;
 wire \data_array.data0[3][42] ;
 wire \data_array.data0[3][43] ;
 wire \data_array.data0[3][44] ;
 wire \data_array.data0[3][45] ;
 wire \data_array.data0[3][46] ;
 wire \data_array.data0[3][47] ;
 wire \data_array.data0[3][48] ;
 wire \data_array.data0[3][49] ;
 wire \data_array.data0[3][4] ;
 wire \data_array.data0[3][50] ;
 wire \data_array.data0[3][51] ;
 wire \data_array.data0[3][52] ;
 wire \data_array.data0[3][53] ;
 wire \data_array.data0[3][54] ;
 wire \data_array.data0[3][55] ;
 wire \data_array.data0[3][56] ;
 wire \data_array.data0[3][57] ;
 wire \data_array.data0[3][58] ;
 wire \data_array.data0[3][59] ;
 wire \data_array.data0[3][5] ;
 wire \data_array.data0[3][60] ;
 wire \data_array.data0[3][61] ;
 wire \data_array.data0[3][62] ;
 wire \data_array.data0[3][63] ;
 wire \data_array.data0[3][6] ;
 wire \data_array.data0[3][7] ;
 wire \data_array.data0[3][8] ;
 wire \data_array.data0[3][9] ;
 wire \data_array.data0[4][0] ;
 wire \data_array.data0[4][10] ;
 wire \data_array.data0[4][11] ;
 wire \data_array.data0[4][12] ;
 wire \data_array.data0[4][13] ;
 wire \data_array.data0[4][14] ;
 wire \data_array.data0[4][15] ;
 wire \data_array.data0[4][16] ;
 wire \data_array.data0[4][17] ;
 wire \data_array.data0[4][18] ;
 wire \data_array.data0[4][19] ;
 wire \data_array.data0[4][1] ;
 wire \data_array.data0[4][20] ;
 wire \data_array.data0[4][21] ;
 wire \data_array.data0[4][22] ;
 wire \data_array.data0[4][23] ;
 wire \data_array.data0[4][24] ;
 wire \data_array.data0[4][25] ;
 wire \data_array.data0[4][26] ;
 wire \data_array.data0[4][27] ;
 wire \data_array.data0[4][28] ;
 wire \data_array.data0[4][29] ;
 wire \data_array.data0[4][2] ;
 wire \data_array.data0[4][30] ;
 wire \data_array.data0[4][31] ;
 wire \data_array.data0[4][32] ;
 wire \data_array.data0[4][33] ;
 wire \data_array.data0[4][34] ;
 wire \data_array.data0[4][35] ;
 wire \data_array.data0[4][36] ;
 wire \data_array.data0[4][37] ;
 wire \data_array.data0[4][38] ;
 wire \data_array.data0[4][39] ;
 wire \data_array.data0[4][3] ;
 wire \data_array.data0[4][40] ;
 wire \data_array.data0[4][41] ;
 wire \data_array.data0[4][42] ;
 wire \data_array.data0[4][43] ;
 wire \data_array.data0[4][44] ;
 wire \data_array.data0[4][45] ;
 wire \data_array.data0[4][46] ;
 wire \data_array.data0[4][47] ;
 wire \data_array.data0[4][48] ;
 wire \data_array.data0[4][49] ;
 wire \data_array.data0[4][4] ;
 wire \data_array.data0[4][50] ;
 wire \data_array.data0[4][51] ;
 wire \data_array.data0[4][52] ;
 wire \data_array.data0[4][53] ;
 wire \data_array.data0[4][54] ;
 wire \data_array.data0[4][55] ;
 wire \data_array.data0[4][56] ;
 wire \data_array.data0[4][57] ;
 wire \data_array.data0[4][58] ;
 wire \data_array.data0[4][59] ;
 wire \data_array.data0[4][5] ;
 wire \data_array.data0[4][60] ;
 wire \data_array.data0[4][61] ;
 wire \data_array.data0[4][62] ;
 wire \data_array.data0[4][63] ;
 wire \data_array.data0[4][6] ;
 wire \data_array.data0[4][7] ;
 wire \data_array.data0[4][8] ;
 wire \data_array.data0[4][9] ;
 wire \data_array.data0[5][0] ;
 wire \data_array.data0[5][10] ;
 wire \data_array.data0[5][11] ;
 wire \data_array.data0[5][12] ;
 wire \data_array.data0[5][13] ;
 wire \data_array.data0[5][14] ;
 wire \data_array.data0[5][15] ;
 wire \data_array.data0[5][16] ;
 wire \data_array.data0[5][17] ;
 wire \data_array.data0[5][18] ;
 wire \data_array.data0[5][19] ;
 wire \data_array.data0[5][1] ;
 wire \data_array.data0[5][20] ;
 wire \data_array.data0[5][21] ;
 wire \data_array.data0[5][22] ;
 wire \data_array.data0[5][23] ;
 wire \data_array.data0[5][24] ;
 wire \data_array.data0[5][25] ;
 wire \data_array.data0[5][26] ;
 wire \data_array.data0[5][27] ;
 wire \data_array.data0[5][28] ;
 wire \data_array.data0[5][29] ;
 wire \data_array.data0[5][2] ;
 wire \data_array.data0[5][30] ;
 wire \data_array.data0[5][31] ;
 wire \data_array.data0[5][32] ;
 wire \data_array.data0[5][33] ;
 wire \data_array.data0[5][34] ;
 wire \data_array.data0[5][35] ;
 wire \data_array.data0[5][36] ;
 wire \data_array.data0[5][37] ;
 wire \data_array.data0[5][38] ;
 wire \data_array.data0[5][39] ;
 wire \data_array.data0[5][3] ;
 wire \data_array.data0[5][40] ;
 wire \data_array.data0[5][41] ;
 wire \data_array.data0[5][42] ;
 wire \data_array.data0[5][43] ;
 wire \data_array.data0[5][44] ;
 wire \data_array.data0[5][45] ;
 wire \data_array.data0[5][46] ;
 wire \data_array.data0[5][47] ;
 wire \data_array.data0[5][48] ;
 wire \data_array.data0[5][49] ;
 wire \data_array.data0[5][4] ;
 wire \data_array.data0[5][50] ;
 wire \data_array.data0[5][51] ;
 wire \data_array.data0[5][52] ;
 wire \data_array.data0[5][53] ;
 wire \data_array.data0[5][54] ;
 wire \data_array.data0[5][55] ;
 wire \data_array.data0[5][56] ;
 wire \data_array.data0[5][57] ;
 wire \data_array.data0[5][58] ;
 wire \data_array.data0[5][59] ;
 wire \data_array.data0[5][5] ;
 wire \data_array.data0[5][60] ;
 wire \data_array.data0[5][61] ;
 wire \data_array.data0[5][62] ;
 wire \data_array.data0[5][63] ;
 wire \data_array.data0[5][6] ;
 wire \data_array.data0[5][7] ;
 wire \data_array.data0[5][8] ;
 wire \data_array.data0[5][9] ;
 wire \data_array.data0[6][0] ;
 wire \data_array.data0[6][10] ;
 wire \data_array.data0[6][11] ;
 wire \data_array.data0[6][12] ;
 wire \data_array.data0[6][13] ;
 wire \data_array.data0[6][14] ;
 wire \data_array.data0[6][15] ;
 wire \data_array.data0[6][16] ;
 wire \data_array.data0[6][17] ;
 wire \data_array.data0[6][18] ;
 wire \data_array.data0[6][19] ;
 wire \data_array.data0[6][1] ;
 wire \data_array.data0[6][20] ;
 wire \data_array.data0[6][21] ;
 wire \data_array.data0[6][22] ;
 wire \data_array.data0[6][23] ;
 wire \data_array.data0[6][24] ;
 wire \data_array.data0[6][25] ;
 wire \data_array.data0[6][26] ;
 wire \data_array.data0[6][27] ;
 wire \data_array.data0[6][28] ;
 wire \data_array.data0[6][29] ;
 wire \data_array.data0[6][2] ;
 wire \data_array.data0[6][30] ;
 wire \data_array.data0[6][31] ;
 wire \data_array.data0[6][32] ;
 wire \data_array.data0[6][33] ;
 wire \data_array.data0[6][34] ;
 wire \data_array.data0[6][35] ;
 wire \data_array.data0[6][36] ;
 wire \data_array.data0[6][37] ;
 wire \data_array.data0[6][38] ;
 wire \data_array.data0[6][39] ;
 wire \data_array.data0[6][3] ;
 wire \data_array.data0[6][40] ;
 wire \data_array.data0[6][41] ;
 wire \data_array.data0[6][42] ;
 wire \data_array.data0[6][43] ;
 wire \data_array.data0[6][44] ;
 wire \data_array.data0[6][45] ;
 wire \data_array.data0[6][46] ;
 wire \data_array.data0[6][47] ;
 wire \data_array.data0[6][48] ;
 wire \data_array.data0[6][49] ;
 wire \data_array.data0[6][4] ;
 wire \data_array.data0[6][50] ;
 wire \data_array.data0[6][51] ;
 wire \data_array.data0[6][52] ;
 wire \data_array.data0[6][53] ;
 wire \data_array.data0[6][54] ;
 wire \data_array.data0[6][55] ;
 wire \data_array.data0[6][56] ;
 wire \data_array.data0[6][57] ;
 wire \data_array.data0[6][58] ;
 wire \data_array.data0[6][59] ;
 wire \data_array.data0[6][5] ;
 wire \data_array.data0[6][60] ;
 wire \data_array.data0[6][61] ;
 wire \data_array.data0[6][62] ;
 wire \data_array.data0[6][63] ;
 wire \data_array.data0[6][6] ;
 wire \data_array.data0[6][7] ;
 wire \data_array.data0[6][8] ;
 wire \data_array.data0[6][9] ;
 wire \data_array.data0[7][0] ;
 wire \data_array.data0[7][10] ;
 wire \data_array.data0[7][11] ;
 wire \data_array.data0[7][12] ;
 wire \data_array.data0[7][13] ;
 wire \data_array.data0[7][14] ;
 wire \data_array.data0[7][15] ;
 wire \data_array.data0[7][16] ;
 wire \data_array.data0[7][17] ;
 wire \data_array.data0[7][18] ;
 wire \data_array.data0[7][19] ;
 wire \data_array.data0[7][1] ;
 wire \data_array.data0[7][20] ;
 wire \data_array.data0[7][21] ;
 wire \data_array.data0[7][22] ;
 wire \data_array.data0[7][23] ;
 wire \data_array.data0[7][24] ;
 wire \data_array.data0[7][25] ;
 wire \data_array.data0[7][26] ;
 wire \data_array.data0[7][27] ;
 wire \data_array.data0[7][28] ;
 wire \data_array.data0[7][29] ;
 wire \data_array.data0[7][2] ;
 wire \data_array.data0[7][30] ;
 wire \data_array.data0[7][31] ;
 wire \data_array.data0[7][32] ;
 wire \data_array.data0[7][33] ;
 wire \data_array.data0[7][34] ;
 wire \data_array.data0[7][35] ;
 wire \data_array.data0[7][36] ;
 wire \data_array.data0[7][37] ;
 wire \data_array.data0[7][38] ;
 wire \data_array.data0[7][39] ;
 wire \data_array.data0[7][3] ;
 wire \data_array.data0[7][40] ;
 wire \data_array.data0[7][41] ;
 wire \data_array.data0[7][42] ;
 wire \data_array.data0[7][43] ;
 wire \data_array.data0[7][44] ;
 wire \data_array.data0[7][45] ;
 wire \data_array.data0[7][46] ;
 wire \data_array.data0[7][47] ;
 wire \data_array.data0[7][48] ;
 wire \data_array.data0[7][49] ;
 wire \data_array.data0[7][4] ;
 wire \data_array.data0[7][50] ;
 wire \data_array.data0[7][51] ;
 wire \data_array.data0[7][52] ;
 wire \data_array.data0[7][53] ;
 wire \data_array.data0[7][54] ;
 wire \data_array.data0[7][55] ;
 wire \data_array.data0[7][56] ;
 wire \data_array.data0[7][57] ;
 wire \data_array.data0[7][58] ;
 wire \data_array.data0[7][59] ;
 wire \data_array.data0[7][5] ;
 wire \data_array.data0[7][60] ;
 wire \data_array.data0[7][61] ;
 wire \data_array.data0[7][62] ;
 wire \data_array.data0[7][63] ;
 wire \data_array.data0[7][6] ;
 wire \data_array.data0[7][7] ;
 wire \data_array.data0[7][8] ;
 wire \data_array.data0[7][9] ;
 wire \data_array.data0[8][0] ;
 wire \data_array.data0[8][10] ;
 wire \data_array.data0[8][11] ;
 wire \data_array.data0[8][12] ;
 wire \data_array.data0[8][13] ;
 wire \data_array.data0[8][14] ;
 wire \data_array.data0[8][15] ;
 wire \data_array.data0[8][16] ;
 wire \data_array.data0[8][17] ;
 wire \data_array.data0[8][18] ;
 wire \data_array.data0[8][19] ;
 wire \data_array.data0[8][1] ;
 wire \data_array.data0[8][20] ;
 wire \data_array.data0[8][21] ;
 wire \data_array.data0[8][22] ;
 wire \data_array.data0[8][23] ;
 wire \data_array.data0[8][24] ;
 wire \data_array.data0[8][25] ;
 wire \data_array.data0[8][26] ;
 wire \data_array.data0[8][27] ;
 wire \data_array.data0[8][28] ;
 wire \data_array.data0[8][29] ;
 wire \data_array.data0[8][2] ;
 wire \data_array.data0[8][30] ;
 wire \data_array.data0[8][31] ;
 wire \data_array.data0[8][32] ;
 wire \data_array.data0[8][33] ;
 wire \data_array.data0[8][34] ;
 wire \data_array.data0[8][35] ;
 wire \data_array.data0[8][36] ;
 wire \data_array.data0[8][37] ;
 wire \data_array.data0[8][38] ;
 wire \data_array.data0[8][39] ;
 wire \data_array.data0[8][3] ;
 wire \data_array.data0[8][40] ;
 wire \data_array.data0[8][41] ;
 wire \data_array.data0[8][42] ;
 wire \data_array.data0[8][43] ;
 wire \data_array.data0[8][44] ;
 wire \data_array.data0[8][45] ;
 wire \data_array.data0[8][46] ;
 wire \data_array.data0[8][47] ;
 wire \data_array.data0[8][48] ;
 wire \data_array.data0[8][49] ;
 wire \data_array.data0[8][4] ;
 wire \data_array.data0[8][50] ;
 wire \data_array.data0[8][51] ;
 wire \data_array.data0[8][52] ;
 wire \data_array.data0[8][53] ;
 wire \data_array.data0[8][54] ;
 wire \data_array.data0[8][55] ;
 wire \data_array.data0[8][56] ;
 wire \data_array.data0[8][57] ;
 wire \data_array.data0[8][58] ;
 wire \data_array.data0[8][59] ;
 wire \data_array.data0[8][5] ;
 wire \data_array.data0[8][60] ;
 wire \data_array.data0[8][61] ;
 wire \data_array.data0[8][62] ;
 wire \data_array.data0[8][63] ;
 wire \data_array.data0[8][6] ;
 wire \data_array.data0[8][7] ;
 wire \data_array.data0[8][8] ;
 wire \data_array.data0[8][9] ;
 wire \data_array.data0[9][0] ;
 wire \data_array.data0[9][10] ;
 wire \data_array.data0[9][11] ;
 wire \data_array.data0[9][12] ;
 wire \data_array.data0[9][13] ;
 wire \data_array.data0[9][14] ;
 wire \data_array.data0[9][15] ;
 wire \data_array.data0[9][16] ;
 wire \data_array.data0[9][17] ;
 wire \data_array.data0[9][18] ;
 wire \data_array.data0[9][19] ;
 wire \data_array.data0[9][1] ;
 wire \data_array.data0[9][20] ;
 wire \data_array.data0[9][21] ;
 wire \data_array.data0[9][22] ;
 wire \data_array.data0[9][23] ;
 wire \data_array.data0[9][24] ;
 wire \data_array.data0[9][25] ;
 wire \data_array.data0[9][26] ;
 wire \data_array.data0[9][27] ;
 wire \data_array.data0[9][28] ;
 wire \data_array.data0[9][29] ;
 wire \data_array.data0[9][2] ;
 wire \data_array.data0[9][30] ;
 wire \data_array.data0[9][31] ;
 wire \data_array.data0[9][32] ;
 wire \data_array.data0[9][33] ;
 wire \data_array.data0[9][34] ;
 wire \data_array.data0[9][35] ;
 wire \data_array.data0[9][36] ;
 wire \data_array.data0[9][37] ;
 wire \data_array.data0[9][38] ;
 wire \data_array.data0[9][39] ;
 wire \data_array.data0[9][3] ;
 wire \data_array.data0[9][40] ;
 wire \data_array.data0[9][41] ;
 wire \data_array.data0[9][42] ;
 wire \data_array.data0[9][43] ;
 wire \data_array.data0[9][44] ;
 wire \data_array.data0[9][45] ;
 wire \data_array.data0[9][46] ;
 wire \data_array.data0[9][47] ;
 wire \data_array.data0[9][48] ;
 wire \data_array.data0[9][49] ;
 wire \data_array.data0[9][4] ;
 wire \data_array.data0[9][50] ;
 wire \data_array.data0[9][51] ;
 wire \data_array.data0[9][52] ;
 wire \data_array.data0[9][53] ;
 wire \data_array.data0[9][54] ;
 wire \data_array.data0[9][55] ;
 wire \data_array.data0[9][56] ;
 wire \data_array.data0[9][57] ;
 wire \data_array.data0[9][58] ;
 wire \data_array.data0[9][59] ;
 wire \data_array.data0[9][5] ;
 wire \data_array.data0[9][60] ;
 wire \data_array.data0[9][61] ;
 wire \data_array.data0[9][62] ;
 wire \data_array.data0[9][63] ;
 wire \data_array.data0[9][6] ;
 wire \data_array.data0[9][7] ;
 wire \data_array.data0[9][8] ;
 wire \data_array.data0[9][9] ;
 wire \data_array.data1[0][0] ;
 wire \data_array.data1[0][10] ;
 wire \data_array.data1[0][11] ;
 wire \data_array.data1[0][12] ;
 wire \data_array.data1[0][13] ;
 wire \data_array.data1[0][14] ;
 wire \data_array.data1[0][15] ;
 wire \data_array.data1[0][16] ;
 wire \data_array.data1[0][17] ;
 wire \data_array.data1[0][18] ;
 wire \data_array.data1[0][19] ;
 wire \data_array.data1[0][1] ;
 wire \data_array.data1[0][20] ;
 wire \data_array.data1[0][21] ;
 wire \data_array.data1[0][22] ;
 wire \data_array.data1[0][23] ;
 wire \data_array.data1[0][24] ;
 wire \data_array.data1[0][25] ;
 wire \data_array.data1[0][26] ;
 wire \data_array.data1[0][27] ;
 wire \data_array.data1[0][28] ;
 wire \data_array.data1[0][29] ;
 wire \data_array.data1[0][2] ;
 wire \data_array.data1[0][30] ;
 wire \data_array.data1[0][31] ;
 wire \data_array.data1[0][32] ;
 wire \data_array.data1[0][33] ;
 wire \data_array.data1[0][34] ;
 wire \data_array.data1[0][35] ;
 wire \data_array.data1[0][36] ;
 wire \data_array.data1[0][37] ;
 wire \data_array.data1[0][38] ;
 wire \data_array.data1[0][39] ;
 wire \data_array.data1[0][3] ;
 wire \data_array.data1[0][40] ;
 wire \data_array.data1[0][41] ;
 wire \data_array.data1[0][42] ;
 wire \data_array.data1[0][43] ;
 wire \data_array.data1[0][44] ;
 wire \data_array.data1[0][45] ;
 wire \data_array.data1[0][46] ;
 wire \data_array.data1[0][47] ;
 wire \data_array.data1[0][48] ;
 wire \data_array.data1[0][49] ;
 wire \data_array.data1[0][4] ;
 wire \data_array.data1[0][50] ;
 wire \data_array.data1[0][51] ;
 wire \data_array.data1[0][52] ;
 wire \data_array.data1[0][53] ;
 wire \data_array.data1[0][54] ;
 wire \data_array.data1[0][55] ;
 wire \data_array.data1[0][56] ;
 wire \data_array.data1[0][57] ;
 wire \data_array.data1[0][58] ;
 wire \data_array.data1[0][59] ;
 wire \data_array.data1[0][5] ;
 wire \data_array.data1[0][60] ;
 wire \data_array.data1[0][61] ;
 wire \data_array.data1[0][62] ;
 wire \data_array.data1[0][63] ;
 wire \data_array.data1[0][6] ;
 wire \data_array.data1[0][7] ;
 wire \data_array.data1[0][8] ;
 wire \data_array.data1[0][9] ;
 wire \data_array.data1[10][0] ;
 wire \data_array.data1[10][10] ;
 wire \data_array.data1[10][11] ;
 wire \data_array.data1[10][12] ;
 wire \data_array.data1[10][13] ;
 wire \data_array.data1[10][14] ;
 wire \data_array.data1[10][15] ;
 wire \data_array.data1[10][16] ;
 wire \data_array.data1[10][17] ;
 wire \data_array.data1[10][18] ;
 wire \data_array.data1[10][19] ;
 wire \data_array.data1[10][1] ;
 wire \data_array.data1[10][20] ;
 wire \data_array.data1[10][21] ;
 wire \data_array.data1[10][22] ;
 wire \data_array.data1[10][23] ;
 wire \data_array.data1[10][24] ;
 wire \data_array.data1[10][25] ;
 wire \data_array.data1[10][26] ;
 wire \data_array.data1[10][27] ;
 wire \data_array.data1[10][28] ;
 wire \data_array.data1[10][29] ;
 wire \data_array.data1[10][2] ;
 wire \data_array.data1[10][30] ;
 wire \data_array.data1[10][31] ;
 wire \data_array.data1[10][32] ;
 wire \data_array.data1[10][33] ;
 wire \data_array.data1[10][34] ;
 wire \data_array.data1[10][35] ;
 wire \data_array.data1[10][36] ;
 wire \data_array.data1[10][37] ;
 wire \data_array.data1[10][38] ;
 wire \data_array.data1[10][39] ;
 wire \data_array.data1[10][3] ;
 wire \data_array.data1[10][40] ;
 wire \data_array.data1[10][41] ;
 wire \data_array.data1[10][42] ;
 wire \data_array.data1[10][43] ;
 wire \data_array.data1[10][44] ;
 wire \data_array.data1[10][45] ;
 wire \data_array.data1[10][46] ;
 wire \data_array.data1[10][47] ;
 wire \data_array.data1[10][48] ;
 wire \data_array.data1[10][49] ;
 wire \data_array.data1[10][4] ;
 wire \data_array.data1[10][50] ;
 wire \data_array.data1[10][51] ;
 wire \data_array.data1[10][52] ;
 wire \data_array.data1[10][53] ;
 wire \data_array.data1[10][54] ;
 wire \data_array.data1[10][55] ;
 wire \data_array.data1[10][56] ;
 wire \data_array.data1[10][57] ;
 wire \data_array.data1[10][58] ;
 wire \data_array.data1[10][59] ;
 wire \data_array.data1[10][5] ;
 wire \data_array.data1[10][60] ;
 wire \data_array.data1[10][61] ;
 wire \data_array.data1[10][62] ;
 wire \data_array.data1[10][63] ;
 wire \data_array.data1[10][6] ;
 wire \data_array.data1[10][7] ;
 wire \data_array.data1[10][8] ;
 wire \data_array.data1[10][9] ;
 wire \data_array.data1[11][0] ;
 wire \data_array.data1[11][10] ;
 wire \data_array.data1[11][11] ;
 wire \data_array.data1[11][12] ;
 wire \data_array.data1[11][13] ;
 wire \data_array.data1[11][14] ;
 wire \data_array.data1[11][15] ;
 wire \data_array.data1[11][16] ;
 wire \data_array.data1[11][17] ;
 wire \data_array.data1[11][18] ;
 wire \data_array.data1[11][19] ;
 wire \data_array.data1[11][1] ;
 wire \data_array.data1[11][20] ;
 wire \data_array.data1[11][21] ;
 wire \data_array.data1[11][22] ;
 wire \data_array.data1[11][23] ;
 wire \data_array.data1[11][24] ;
 wire \data_array.data1[11][25] ;
 wire \data_array.data1[11][26] ;
 wire \data_array.data1[11][27] ;
 wire \data_array.data1[11][28] ;
 wire \data_array.data1[11][29] ;
 wire \data_array.data1[11][2] ;
 wire \data_array.data1[11][30] ;
 wire \data_array.data1[11][31] ;
 wire \data_array.data1[11][32] ;
 wire \data_array.data1[11][33] ;
 wire \data_array.data1[11][34] ;
 wire \data_array.data1[11][35] ;
 wire \data_array.data1[11][36] ;
 wire \data_array.data1[11][37] ;
 wire \data_array.data1[11][38] ;
 wire \data_array.data1[11][39] ;
 wire \data_array.data1[11][3] ;
 wire \data_array.data1[11][40] ;
 wire \data_array.data1[11][41] ;
 wire \data_array.data1[11][42] ;
 wire \data_array.data1[11][43] ;
 wire \data_array.data1[11][44] ;
 wire \data_array.data1[11][45] ;
 wire \data_array.data1[11][46] ;
 wire \data_array.data1[11][47] ;
 wire \data_array.data1[11][48] ;
 wire \data_array.data1[11][49] ;
 wire \data_array.data1[11][4] ;
 wire \data_array.data1[11][50] ;
 wire \data_array.data1[11][51] ;
 wire \data_array.data1[11][52] ;
 wire \data_array.data1[11][53] ;
 wire \data_array.data1[11][54] ;
 wire \data_array.data1[11][55] ;
 wire \data_array.data1[11][56] ;
 wire \data_array.data1[11][57] ;
 wire \data_array.data1[11][58] ;
 wire \data_array.data1[11][59] ;
 wire \data_array.data1[11][5] ;
 wire \data_array.data1[11][60] ;
 wire \data_array.data1[11][61] ;
 wire \data_array.data1[11][62] ;
 wire \data_array.data1[11][63] ;
 wire \data_array.data1[11][6] ;
 wire \data_array.data1[11][7] ;
 wire \data_array.data1[11][8] ;
 wire \data_array.data1[11][9] ;
 wire \data_array.data1[12][0] ;
 wire \data_array.data1[12][10] ;
 wire \data_array.data1[12][11] ;
 wire \data_array.data1[12][12] ;
 wire \data_array.data1[12][13] ;
 wire \data_array.data1[12][14] ;
 wire \data_array.data1[12][15] ;
 wire \data_array.data1[12][16] ;
 wire \data_array.data1[12][17] ;
 wire \data_array.data1[12][18] ;
 wire \data_array.data1[12][19] ;
 wire \data_array.data1[12][1] ;
 wire \data_array.data1[12][20] ;
 wire \data_array.data1[12][21] ;
 wire \data_array.data1[12][22] ;
 wire \data_array.data1[12][23] ;
 wire \data_array.data1[12][24] ;
 wire \data_array.data1[12][25] ;
 wire \data_array.data1[12][26] ;
 wire \data_array.data1[12][27] ;
 wire \data_array.data1[12][28] ;
 wire \data_array.data1[12][29] ;
 wire \data_array.data1[12][2] ;
 wire \data_array.data1[12][30] ;
 wire \data_array.data1[12][31] ;
 wire \data_array.data1[12][32] ;
 wire \data_array.data1[12][33] ;
 wire \data_array.data1[12][34] ;
 wire \data_array.data1[12][35] ;
 wire \data_array.data1[12][36] ;
 wire \data_array.data1[12][37] ;
 wire \data_array.data1[12][38] ;
 wire \data_array.data1[12][39] ;
 wire \data_array.data1[12][3] ;
 wire \data_array.data1[12][40] ;
 wire \data_array.data1[12][41] ;
 wire \data_array.data1[12][42] ;
 wire \data_array.data1[12][43] ;
 wire \data_array.data1[12][44] ;
 wire \data_array.data1[12][45] ;
 wire \data_array.data1[12][46] ;
 wire \data_array.data1[12][47] ;
 wire \data_array.data1[12][48] ;
 wire \data_array.data1[12][49] ;
 wire \data_array.data1[12][4] ;
 wire \data_array.data1[12][50] ;
 wire \data_array.data1[12][51] ;
 wire \data_array.data1[12][52] ;
 wire \data_array.data1[12][53] ;
 wire \data_array.data1[12][54] ;
 wire \data_array.data1[12][55] ;
 wire \data_array.data1[12][56] ;
 wire \data_array.data1[12][57] ;
 wire \data_array.data1[12][58] ;
 wire \data_array.data1[12][59] ;
 wire \data_array.data1[12][5] ;
 wire \data_array.data1[12][60] ;
 wire \data_array.data1[12][61] ;
 wire \data_array.data1[12][62] ;
 wire \data_array.data1[12][63] ;
 wire \data_array.data1[12][6] ;
 wire \data_array.data1[12][7] ;
 wire \data_array.data1[12][8] ;
 wire \data_array.data1[12][9] ;
 wire \data_array.data1[13][0] ;
 wire \data_array.data1[13][10] ;
 wire \data_array.data1[13][11] ;
 wire \data_array.data1[13][12] ;
 wire \data_array.data1[13][13] ;
 wire \data_array.data1[13][14] ;
 wire \data_array.data1[13][15] ;
 wire \data_array.data1[13][16] ;
 wire \data_array.data1[13][17] ;
 wire \data_array.data1[13][18] ;
 wire \data_array.data1[13][19] ;
 wire \data_array.data1[13][1] ;
 wire \data_array.data1[13][20] ;
 wire \data_array.data1[13][21] ;
 wire \data_array.data1[13][22] ;
 wire \data_array.data1[13][23] ;
 wire \data_array.data1[13][24] ;
 wire \data_array.data1[13][25] ;
 wire \data_array.data1[13][26] ;
 wire \data_array.data1[13][27] ;
 wire \data_array.data1[13][28] ;
 wire \data_array.data1[13][29] ;
 wire \data_array.data1[13][2] ;
 wire \data_array.data1[13][30] ;
 wire \data_array.data1[13][31] ;
 wire \data_array.data1[13][32] ;
 wire \data_array.data1[13][33] ;
 wire \data_array.data1[13][34] ;
 wire \data_array.data1[13][35] ;
 wire \data_array.data1[13][36] ;
 wire \data_array.data1[13][37] ;
 wire \data_array.data1[13][38] ;
 wire \data_array.data1[13][39] ;
 wire \data_array.data1[13][3] ;
 wire \data_array.data1[13][40] ;
 wire \data_array.data1[13][41] ;
 wire \data_array.data1[13][42] ;
 wire \data_array.data1[13][43] ;
 wire \data_array.data1[13][44] ;
 wire \data_array.data1[13][45] ;
 wire \data_array.data1[13][46] ;
 wire \data_array.data1[13][47] ;
 wire \data_array.data1[13][48] ;
 wire \data_array.data1[13][49] ;
 wire \data_array.data1[13][4] ;
 wire \data_array.data1[13][50] ;
 wire \data_array.data1[13][51] ;
 wire \data_array.data1[13][52] ;
 wire \data_array.data1[13][53] ;
 wire \data_array.data1[13][54] ;
 wire \data_array.data1[13][55] ;
 wire \data_array.data1[13][56] ;
 wire \data_array.data1[13][57] ;
 wire \data_array.data1[13][58] ;
 wire \data_array.data1[13][59] ;
 wire \data_array.data1[13][5] ;
 wire \data_array.data1[13][60] ;
 wire \data_array.data1[13][61] ;
 wire \data_array.data1[13][62] ;
 wire \data_array.data1[13][63] ;
 wire \data_array.data1[13][6] ;
 wire \data_array.data1[13][7] ;
 wire \data_array.data1[13][8] ;
 wire \data_array.data1[13][9] ;
 wire \data_array.data1[14][0] ;
 wire \data_array.data1[14][10] ;
 wire \data_array.data1[14][11] ;
 wire \data_array.data1[14][12] ;
 wire \data_array.data1[14][13] ;
 wire \data_array.data1[14][14] ;
 wire \data_array.data1[14][15] ;
 wire \data_array.data1[14][16] ;
 wire \data_array.data1[14][17] ;
 wire \data_array.data1[14][18] ;
 wire \data_array.data1[14][19] ;
 wire \data_array.data1[14][1] ;
 wire \data_array.data1[14][20] ;
 wire \data_array.data1[14][21] ;
 wire \data_array.data1[14][22] ;
 wire \data_array.data1[14][23] ;
 wire \data_array.data1[14][24] ;
 wire \data_array.data1[14][25] ;
 wire \data_array.data1[14][26] ;
 wire \data_array.data1[14][27] ;
 wire \data_array.data1[14][28] ;
 wire \data_array.data1[14][29] ;
 wire \data_array.data1[14][2] ;
 wire \data_array.data1[14][30] ;
 wire \data_array.data1[14][31] ;
 wire \data_array.data1[14][32] ;
 wire \data_array.data1[14][33] ;
 wire \data_array.data1[14][34] ;
 wire \data_array.data1[14][35] ;
 wire \data_array.data1[14][36] ;
 wire \data_array.data1[14][37] ;
 wire \data_array.data1[14][38] ;
 wire \data_array.data1[14][39] ;
 wire \data_array.data1[14][3] ;
 wire \data_array.data1[14][40] ;
 wire \data_array.data1[14][41] ;
 wire \data_array.data1[14][42] ;
 wire \data_array.data1[14][43] ;
 wire \data_array.data1[14][44] ;
 wire \data_array.data1[14][45] ;
 wire \data_array.data1[14][46] ;
 wire \data_array.data1[14][47] ;
 wire \data_array.data1[14][48] ;
 wire \data_array.data1[14][49] ;
 wire \data_array.data1[14][4] ;
 wire \data_array.data1[14][50] ;
 wire \data_array.data1[14][51] ;
 wire \data_array.data1[14][52] ;
 wire \data_array.data1[14][53] ;
 wire \data_array.data1[14][54] ;
 wire \data_array.data1[14][55] ;
 wire \data_array.data1[14][56] ;
 wire \data_array.data1[14][57] ;
 wire \data_array.data1[14][58] ;
 wire \data_array.data1[14][59] ;
 wire \data_array.data1[14][5] ;
 wire \data_array.data1[14][60] ;
 wire \data_array.data1[14][61] ;
 wire \data_array.data1[14][62] ;
 wire \data_array.data1[14][63] ;
 wire \data_array.data1[14][6] ;
 wire \data_array.data1[14][7] ;
 wire \data_array.data1[14][8] ;
 wire \data_array.data1[14][9] ;
 wire \data_array.data1[15][0] ;
 wire \data_array.data1[15][10] ;
 wire \data_array.data1[15][11] ;
 wire \data_array.data1[15][12] ;
 wire \data_array.data1[15][13] ;
 wire \data_array.data1[15][14] ;
 wire \data_array.data1[15][15] ;
 wire \data_array.data1[15][16] ;
 wire \data_array.data1[15][17] ;
 wire \data_array.data1[15][18] ;
 wire \data_array.data1[15][19] ;
 wire \data_array.data1[15][1] ;
 wire \data_array.data1[15][20] ;
 wire \data_array.data1[15][21] ;
 wire \data_array.data1[15][22] ;
 wire \data_array.data1[15][23] ;
 wire \data_array.data1[15][24] ;
 wire \data_array.data1[15][25] ;
 wire \data_array.data1[15][26] ;
 wire \data_array.data1[15][27] ;
 wire \data_array.data1[15][28] ;
 wire \data_array.data1[15][29] ;
 wire \data_array.data1[15][2] ;
 wire \data_array.data1[15][30] ;
 wire \data_array.data1[15][31] ;
 wire \data_array.data1[15][32] ;
 wire \data_array.data1[15][33] ;
 wire \data_array.data1[15][34] ;
 wire \data_array.data1[15][35] ;
 wire \data_array.data1[15][36] ;
 wire \data_array.data1[15][37] ;
 wire \data_array.data1[15][38] ;
 wire \data_array.data1[15][39] ;
 wire \data_array.data1[15][3] ;
 wire \data_array.data1[15][40] ;
 wire \data_array.data1[15][41] ;
 wire \data_array.data1[15][42] ;
 wire \data_array.data1[15][43] ;
 wire \data_array.data1[15][44] ;
 wire \data_array.data1[15][45] ;
 wire \data_array.data1[15][46] ;
 wire \data_array.data1[15][47] ;
 wire \data_array.data1[15][48] ;
 wire \data_array.data1[15][49] ;
 wire \data_array.data1[15][4] ;
 wire \data_array.data1[15][50] ;
 wire \data_array.data1[15][51] ;
 wire \data_array.data1[15][52] ;
 wire \data_array.data1[15][53] ;
 wire \data_array.data1[15][54] ;
 wire \data_array.data1[15][55] ;
 wire \data_array.data1[15][56] ;
 wire \data_array.data1[15][57] ;
 wire \data_array.data1[15][58] ;
 wire \data_array.data1[15][59] ;
 wire \data_array.data1[15][5] ;
 wire \data_array.data1[15][60] ;
 wire \data_array.data1[15][61] ;
 wire \data_array.data1[15][62] ;
 wire \data_array.data1[15][63] ;
 wire \data_array.data1[15][6] ;
 wire \data_array.data1[15][7] ;
 wire \data_array.data1[15][8] ;
 wire \data_array.data1[15][9] ;
 wire \data_array.data1[1][0] ;
 wire \data_array.data1[1][10] ;
 wire \data_array.data1[1][11] ;
 wire \data_array.data1[1][12] ;
 wire \data_array.data1[1][13] ;
 wire \data_array.data1[1][14] ;
 wire \data_array.data1[1][15] ;
 wire \data_array.data1[1][16] ;
 wire \data_array.data1[1][17] ;
 wire \data_array.data1[1][18] ;
 wire \data_array.data1[1][19] ;
 wire \data_array.data1[1][1] ;
 wire \data_array.data1[1][20] ;
 wire \data_array.data1[1][21] ;
 wire \data_array.data1[1][22] ;
 wire \data_array.data1[1][23] ;
 wire \data_array.data1[1][24] ;
 wire \data_array.data1[1][25] ;
 wire \data_array.data1[1][26] ;
 wire \data_array.data1[1][27] ;
 wire \data_array.data1[1][28] ;
 wire \data_array.data1[1][29] ;
 wire \data_array.data1[1][2] ;
 wire \data_array.data1[1][30] ;
 wire \data_array.data1[1][31] ;
 wire \data_array.data1[1][32] ;
 wire \data_array.data1[1][33] ;
 wire \data_array.data1[1][34] ;
 wire \data_array.data1[1][35] ;
 wire \data_array.data1[1][36] ;
 wire \data_array.data1[1][37] ;
 wire \data_array.data1[1][38] ;
 wire \data_array.data1[1][39] ;
 wire \data_array.data1[1][3] ;
 wire \data_array.data1[1][40] ;
 wire \data_array.data1[1][41] ;
 wire \data_array.data1[1][42] ;
 wire \data_array.data1[1][43] ;
 wire \data_array.data1[1][44] ;
 wire \data_array.data1[1][45] ;
 wire \data_array.data1[1][46] ;
 wire \data_array.data1[1][47] ;
 wire \data_array.data1[1][48] ;
 wire \data_array.data1[1][49] ;
 wire \data_array.data1[1][4] ;
 wire \data_array.data1[1][50] ;
 wire \data_array.data1[1][51] ;
 wire \data_array.data1[1][52] ;
 wire \data_array.data1[1][53] ;
 wire \data_array.data1[1][54] ;
 wire \data_array.data1[1][55] ;
 wire \data_array.data1[1][56] ;
 wire \data_array.data1[1][57] ;
 wire \data_array.data1[1][58] ;
 wire \data_array.data1[1][59] ;
 wire \data_array.data1[1][5] ;
 wire \data_array.data1[1][60] ;
 wire \data_array.data1[1][61] ;
 wire \data_array.data1[1][62] ;
 wire \data_array.data1[1][63] ;
 wire \data_array.data1[1][6] ;
 wire \data_array.data1[1][7] ;
 wire \data_array.data1[1][8] ;
 wire \data_array.data1[1][9] ;
 wire \data_array.data1[2][0] ;
 wire \data_array.data1[2][10] ;
 wire \data_array.data1[2][11] ;
 wire \data_array.data1[2][12] ;
 wire \data_array.data1[2][13] ;
 wire \data_array.data1[2][14] ;
 wire \data_array.data1[2][15] ;
 wire \data_array.data1[2][16] ;
 wire \data_array.data1[2][17] ;
 wire \data_array.data1[2][18] ;
 wire \data_array.data1[2][19] ;
 wire \data_array.data1[2][1] ;
 wire \data_array.data1[2][20] ;
 wire \data_array.data1[2][21] ;
 wire \data_array.data1[2][22] ;
 wire \data_array.data1[2][23] ;
 wire \data_array.data1[2][24] ;
 wire \data_array.data1[2][25] ;
 wire \data_array.data1[2][26] ;
 wire \data_array.data1[2][27] ;
 wire \data_array.data1[2][28] ;
 wire \data_array.data1[2][29] ;
 wire \data_array.data1[2][2] ;
 wire \data_array.data1[2][30] ;
 wire \data_array.data1[2][31] ;
 wire \data_array.data1[2][32] ;
 wire \data_array.data1[2][33] ;
 wire \data_array.data1[2][34] ;
 wire \data_array.data1[2][35] ;
 wire \data_array.data1[2][36] ;
 wire \data_array.data1[2][37] ;
 wire \data_array.data1[2][38] ;
 wire \data_array.data1[2][39] ;
 wire \data_array.data1[2][3] ;
 wire \data_array.data1[2][40] ;
 wire \data_array.data1[2][41] ;
 wire \data_array.data1[2][42] ;
 wire \data_array.data1[2][43] ;
 wire \data_array.data1[2][44] ;
 wire \data_array.data1[2][45] ;
 wire \data_array.data1[2][46] ;
 wire \data_array.data1[2][47] ;
 wire \data_array.data1[2][48] ;
 wire \data_array.data1[2][49] ;
 wire \data_array.data1[2][4] ;
 wire \data_array.data1[2][50] ;
 wire \data_array.data1[2][51] ;
 wire \data_array.data1[2][52] ;
 wire \data_array.data1[2][53] ;
 wire \data_array.data1[2][54] ;
 wire \data_array.data1[2][55] ;
 wire \data_array.data1[2][56] ;
 wire \data_array.data1[2][57] ;
 wire \data_array.data1[2][58] ;
 wire \data_array.data1[2][59] ;
 wire \data_array.data1[2][5] ;
 wire \data_array.data1[2][60] ;
 wire \data_array.data1[2][61] ;
 wire \data_array.data1[2][62] ;
 wire \data_array.data1[2][63] ;
 wire \data_array.data1[2][6] ;
 wire \data_array.data1[2][7] ;
 wire \data_array.data1[2][8] ;
 wire \data_array.data1[2][9] ;
 wire \data_array.data1[3][0] ;
 wire \data_array.data1[3][10] ;
 wire \data_array.data1[3][11] ;
 wire \data_array.data1[3][12] ;
 wire \data_array.data1[3][13] ;
 wire \data_array.data1[3][14] ;
 wire \data_array.data1[3][15] ;
 wire \data_array.data1[3][16] ;
 wire \data_array.data1[3][17] ;
 wire \data_array.data1[3][18] ;
 wire \data_array.data1[3][19] ;
 wire \data_array.data1[3][1] ;
 wire \data_array.data1[3][20] ;
 wire \data_array.data1[3][21] ;
 wire \data_array.data1[3][22] ;
 wire \data_array.data1[3][23] ;
 wire \data_array.data1[3][24] ;
 wire \data_array.data1[3][25] ;
 wire \data_array.data1[3][26] ;
 wire \data_array.data1[3][27] ;
 wire \data_array.data1[3][28] ;
 wire \data_array.data1[3][29] ;
 wire \data_array.data1[3][2] ;
 wire \data_array.data1[3][30] ;
 wire \data_array.data1[3][31] ;
 wire \data_array.data1[3][32] ;
 wire \data_array.data1[3][33] ;
 wire \data_array.data1[3][34] ;
 wire \data_array.data1[3][35] ;
 wire \data_array.data1[3][36] ;
 wire \data_array.data1[3][37] ;
 wire \data_array.data1[3][38] ;
 wire \data_array.data1[3][39] ;
 wire \data_array.data1[3][3] ;
 wire \data_array.data1[3][40] ;
 wire \data_array.data1[3][41] ;
 wire \data_array.data1[3][42] ;
 wire \data_array.data1[3][43] ;
 wire \data_array.data1[3][44] ;
 wire \data_array.data1[3][45] ;
 wire \data_array.data1[3][46] ;
 wire \data_array.data1[3][47] ;
 wire \data_array.data1[3][48] ;
 wire \data_array.data1[3][49] ;
 wire \data_array.data1[3][4] ;
 wire \data_array.data1[3][50] ;
 wire \data_array.data1[3][51] ;
 wire \data_array.data1[3][52] ;
 wire \data_array.data1[3][53] ;
 wire \data_array.data1[3][54] ;
 wire \data_array.data1[3][55] ;
 wire \data_array.data1[3][56] ;
 wire \data_array.data1[3][57] ;
 wire \data_array.data1[3][58] ;
 wire \data_array.data1[3][59] ;
 wire \data_array.data1[3][5] ;
 wire \data_array.data1[3][60] ;
 wire \data_array.data1[3][61] ;
 wire \data_array.data1[3][62] ;
 wire \data_array.data1[3][63] ;
 wire \data_array.data1[3][6] ;
 wire \data_array.data1[3][7] ;
 wire \data_array.data1[3][8] ;
 wire \data_array.data1[3][9] ;
 wire \data_array.data1[4][0] ;
 wire \data_array.data1[4][10] ;
 wire \data_array.data1[4][11] ;
 wire \data_array.data1[4][12] ;
 wire \data_array.data1[4][13] ;
 wire \data_array.data1[4][14] ;
 wire \data_array.data1[4][15] ;
 wire \data_array.data1[4][16] ;
 wire \data_array.data1[4][17] ;
 wire \data_array.data1[4][18] ;
 wire \data_array.data1[4][19] ;
 wire \data_array.data1[4][1] ;
 wire \data_array.data1[4][20] ;
 wire \data_array.data1[4][21] ;
 wire \data_array.data1[4][22] ;
 wire \data_array.data1[4][23] ;
 wire \data_array.data1[4][24] ;
 wire \data_array.data1[4][25] ;
 wire \data_array.data1[4][26] ;
 wire \data_array.data1[4][27] ;
 wire \data_array.data1[4][28] ;
 wire \data_array.data1[4][29] ;
 wire \data_array.data1[4][2] ;
 wire \data_array.data1[4][30] ;
 wire \data_array.data1[4][31] ;
 wire \data_array.data1[4][32] ;
 wire \data_array.data1[4][33] ;
 wire \data_array.data1[4][34] ;
 wire \data_array.data1[4][35] ;
 wire \data_array.data1[4][36] ;
 wire \data_array.data1[4][37] ;
 wire \data_array.data1[4][38] ;
 wire \data_array.data1[4][39] ;
 wire \data_array.data1[4][3] ;
 wire \data_array.data1[4][40] ;
 wire \data_array.data1[4][41] ;
 wire \data_array.data1[4][42] ;
 wire \data_array.data1[4][43] ;
 wire \data_array.data1[4][44] ;
 wire \data_array.data1[4][45] ;
 wire \data_array.data1[4][46] ;
 wire \data_array.data1[4][47] ;
 wire \data_array.data1[4][48] ;
 wire \data_array.data1[4][49] ;
 wire \data_array.data1[4][4] ;
 wire \data_array.data1[4][50] ;
 wire \data_array.data1[4][51] ;
 wire \data_array.data1[4][52] ;
 wire \data_array.data1[4][53] ;
 wire \data_array.data1[4][54] ;
 wire \data_array.data1[4][55] ;
 wire \data_array.data1[4][56] ;
 wire \data_array.data1[4][57] ;
 wire \data_array.data1[4][58] ;
 wire \data_array.data1[4][59] ;
 wire \data_array.data1[4][5] ;
 wire \data_array.data1[4][60] ;
 wire \data_array.data1[4][61] ;
 wire \data_array.data1[4][62] ;
 wire \data_array.data1[4][63] ;
 wire \data_array.data1[4][6] ;
 wire \data_array.data1[4][7] ;
 wire \data_array.data1[4][8] ;
 wire \data_array.data1[4][9] ;
 wire \data_array.data1[5][0] ;
 wire \data_array.data1[5][10] ;
 wire \data_array.data1[5][11] ;
 wire \data_array.data1[5][12] ;
 wire \data_array.data1[5][13] ;
 wire \data_array.data1[5][14] ;
 wire \data_array.data1[5][15] ;
 wire \data_array.data1[5][16] ;
 wire \data_array.data1[5][17] ;
 wire \data_array.data1[5][18] ;
 wire \data_array.data1[5][19] ;
 wire \data_array.data1[5][1] ;
 wire \data_array.data1[5][20] ;
 wire \data_array.data1[5][21] ;
 wire \data_array.data1[5][22] ;
 wire \data_array.data1[5][23] ;
 wire \data_array.data1[5][24] ;
 wire \data_array.data1[5][25] ;
 wire \data_array.data1[5][26] ;
 wire \data_array.data1[5][27] ;
 wire \data_array.data1[5][28] ;
 wire \data_array.data1[5][29] ;
 wire \data_array.data1[5][2] ;
 wire \data_array.data1[5][30] ;
 wire \data_array.data1[5][31] ;
 wire \data_array.data1[5][32] ;
 wire \data_array.data1[5][33] ;
 wire \data_array.data1[5][34] ;
 wire \data_array.data1[5][35] ;
 wire \data_array.data1[5][36] ;
 wire \data_array.data1[5][37] ;
 wire \data_array.data1[5][38] ;
 wire \data_array.data1[5][39] ;
 wire \data_array.data1[5][3] ;
 wire \data_array.data1[5][40] ;
 wire \data_array.data1[5][41] ;
 wire \data_array.data1[5][42] ;
 wire \data_array.data1[5][43] ;
 wire \data_array.data1[5][44] ;
 wire \data_array.data1[5][45] ;
 wire \data_array.data1[5][46] ;
 wire \data_array.data1[5][47] ;
 wire \data_array.data1[5][48] ;
 wire \data_array.data1[5][49] ;
 wire \data_array.data1[5][4] ;
 wire \data_array.data1[5][50] ;
 wire \data_array.data1[5][51] ;
 wire \data_array.data1[5][52] ;
 wire \data_array.data1[5][53] ;
 wire \data_array.data1[5][54] ;
 wire \data_array.data1[5][55] ;
 wire \data_array.data1[5][56] ;
 wire \data_array.data1[5][57] ;
 wire \data_array.data1[5][58] ;
 wire \data_array.data1[5][59] ;
 wire \data_array.data1[5][5] ;
 wire \data_array.data1[5][60] ;
 wire \data_array.data1[5][61] ;
 wire \data_array.data1[5][62] ;
 wire \data_array.data1[5][63] ;
 wire \data_array.data1[5][6] ;
 wire \data_array.data1[5][7] ;
 wire \data_array.data1[5][8] ;
 wire \data_array.data1[5][9] ;
 wire \data_array.data1[6][0] ;
 wire \data_array.data1[6][10] ;
 wire \data_array.data1[6][11] ;
 wire \data_array.data1[6][12] ;
 wire \data_array.data1[6][13] ;
 wire \data_array.data1[6][14] ;
 wire \data_array.data1[6][15] ;
 wire \data_array.data1[6][16] ;
 wire \data_array.data1[6][17] ;
 wire \data_array.data1[6][18] ;
 wire \data_array.data1[6][19] ;
 wire \data_array.data1[6][1] ;
 wire \data_array.data1[6][20] ;
 wire \data_array.data1[6][21] ;
 wire \data_array.data1[6][22] ;
 wire \data_array.data1[6][23] ;
 wire \data_array.data1[6][24] ;
 wire \data_array.data1[6][25] ;
 wire \data_array.data1[6][26] ;
 wire \data_array.data1[6][27] ;
 wire \data_array.data1[6][28] ;
 wire \data_array.data1[6][29] ;
 wire \data_array.data1[6][2] ;
 wire \data_array.data1[6][30] ;
 wire \data_array.data1[6][31] ;
 wire \data_array.data1[6][32] ;
 wire \data_array.data1[6][33] ;
 wire \data_array.data1[6][34] ;
 wire \data_array.data1[6][35] ;
 wire \data_array.data1[6][36] ;
 wire \data_array.data1[6][37] ;
 wire \data_array.data1[6][38] ;
 wire \data_array.data1[6][39] ;
 wire \data_array.data1[6][3] ;
 wire \data_array.data1[6][40] ;
 wire \data_array.data1[6][41] ;
 wire \data_array.data1[6][42] ;
 wire \data_array.data1[6][43] ;
 wire \data_array.data1[6][44] ;
 wire \data_array.data1[6][45] ;
 wire \data_array.data1[6][46] ;
 wire \data_array.data1[6][47] ;
 wire \data_array.data1[6][48] ;
 wire \data_array.data1[6][49] ;
 wire \data_array.data1[6][4] ;
 wire \data_array.data1[6][50] ;
 wire \data_array.data1[6][51] ;
 wire \data_array.data1[6][52] ;
 wire \data_array.data1[6][53] ;
 wire \data_array.data1[6][54] ;
 wire \data_array.data1[6][55] ;
 wire \data_array.data1[6][56] ;
 wire \data_array.data1[6][57] ;
 wire \data_array.data1[6][58] ;
 wire \data_array.data1[6][59] ;
 wire \data_array.data1[6][5] ;
 wire \data_array.data1[6][60] ;
 wire \data_array.data1[6][61] ;
 wire \data_array.data1[6][62] ;
 wire \data_array.data1[6][63] ;
 wire \data_array.data1[6][6] ;
 wire \data_array.data1[6][7] ;
 wire \data_array.data1[6][8] ;
 wire \data_array.data1[6][9] ;
 wire \data_array.data1[7][0] ;
 wire \data_array.data1[7][10] ;
 wire \data_array.data1[7][11] ;
 wire \data_array.data1[7][12] ;
 wire \data_array.data1[7][13] ;
 wire \data_array.data1[7][14] ;
 wire \data_array.data1[7][15] ;
 wire \data_array.data1[7][16] ;
 wire \data_array.data1[7][17] ;
 wire \data_array.data1[7][18] ;
 wire \data_array.data1[7][19] ;
 wire \data_array.data1[7][1] ;
 wire \data_array.data1[7][20] ;
 wire \data_array.data1[7][21] ;
 wire \data_array.data1[7][22] ;
 wire \data_array.data1[7][23] ;
 wire \data_array.data1[7][24] ;
 wire \data_array.data1[7][25] ;
 wire \data_array.data1[7][26] ;
 wire \data_array.data1[7][27] ;
 wire \data_array.data1[7][28] ;
 wire \data_array.data1[7][29] ;
 wire \data_array.data1[7][2] ;
 wire \data_array.data1[7][30] ;
 wire \data_array.data1[7][31] ;
 wire \data_array.data1[7][32] ;
 wire \data_array.data1[7][33] ;
 wire \data_array.data1[7][34] ;
 wire \data_array.data1[7][35] ;
 wire \data_array.data1[7][36] ;
 wire \data_array.data1[7][37] ;
 wire \data_array.data1[7][38] ;
 wire \data_array.data1[7][39] ;
 wire \data_array.data1[7][3] ;
 wire \data_array.data1[7][40] ;
 wire \data_array.data1[7][41] ;
 wire \data_array.data1[7][42] ;
 wire \data_array.data1[7][43] ;
 wire \data_array.data1[7][44] ;
 wire \data_array.data1[7][45] ;
 wire \data_array.data1[7][46] ;
 wire \data_array.data1[7][47] ;
 wire \data_array.data1[7][48] ;
 wire \data_array.data1[7][49] ;
 wire \data_array.data1[7][4] ;
 wire \data_array.data1[7][50] ;
 wire \data_array.data1[7][51] ;
 wire \data_array.data1[7][52] ;
 wire \data_array.data1[7][53] ;
 wire \data_array.data1[7][54] ;
 wire \data_array.data1[7][55] ;
 wire \data_array.data1[7][56] ;
 wire \data_array.data1[7][57] ;
 wire \data_array.data1[7][58] ;
 wire \data_array.data1[7][59] ;
 wire \data_array.data1[7][5] ;
 wire \data_array.data1[7][60] ;
 wire \data_array.data1[7][61] ;
 wire \data_array.data1[7][62] ;
 wire \data_array.data1[7][63] ;
 wire \data_array.data1[7][6] ;
 wire \data_array.data1[7][7] ;
 wire \data_array.data1[7][8] ;
 wire \data_array.data1[7][9] ;
 wire \data_array.data1[8][0] ;
 wire \data_array.data1[8][10] ;
 wire \data_array.data1[8][11] ;
 wire \data_array.data1[8][12] ;
 wire \data_array.data1[8][13] ;
 wire \data_array.data1[8][14] ;
 wire \data_array.data1[8][15] ;
 wire \data_array.data1[8][16] ;
 wire \data_array.data1[8][17] ;
 wire \data_array.data1[8][18] ;
 wire \data_array.data1[8][19] ;
 wire \data_array.data1[8][1] ;
 wire \data_array.data1[8][20] ;
 wire \data_array.data1[8][21] ;
 wire \data_array.data1[8][22] ;
 wire \data_array.data1[8][23] ;
 wire \data_array.data1[8][24] ;
 wire \data_array.data1[8][25] ;
 wire \data_array.data1[8][26] ;
 wire \data_array.data1[8][27] ;
 wire \data_array.data1[8][28] ;
 wire \data_array.data1[8][29] ;
 wire \data_array.data1[8][2] ;
 wire \data_array.data1[8][30] ;
 wire \data_array.data1[8][31] ;
 wire \data_array.data1[8][32] ;
 wire \data_array.data1[8][33] ;
 wire \data_array.data1[8][34] ;
 wire \data_array.data1[8][35] ;
 wire \data_array.data1[8][36] ;
 wire \data_array.data1[8][37] ;
 wire \data_array.data1[8][38] ;
 wire \data_array.data1[8][39] ;
 wire \data_array.data1[8][3] ;
 wire \data_array.data1[8][40] ;
 wire \data_array.data1[8][41] ;
 wire \data_array.data1[8][42] ;
 wire \data_array.data1[8][43] ;
 wire \data_array.data1[8][44] ;
 wire \data_array.data1[8][45] ;
 wire \data_array.data1[8][46] ;
 wire \data_array.data1[8][47] ;
 wire \data_array.data1[8][48] ;
 wire \data_array.data1[8][49] ;
 wire \data_array.data1[8][4] ;
 wire \data_array.data1[8][50] ;
 wire \data_array.data1[8][51] ;
 wire \data_array.data1[8][52] ;
 wire \data_array.data1[8][53] ;
 wire \data_array.data1[8][54] ;
 wire \data_array.data1[8][55] ;
 wire \data_array.data1[8][56] ;
 wire \data_array.data1[8][57] ;
 wire \data_array.data1[8][58] ;
 wire \data_array.data1[8][59] ;
 wire \data_array.data1[8][5] ;
 wire \data_array.data1[8][60] ;
 wire \data_array.data1[8][61] ;
 wire \data_array.data1[8][62] ;
 wire \data_array.data1[8][63] ;
 wire \data_array.data1[8][6] ;
 wire \data_array.data1[8][7] ;
 wire \data_array.data1[8][8] ;
 wire \data_array.data1[8][9] ;
 wire \data_array.data1[9][0] ;
 wire \data_array.data1[9][10] ;
 wire \data_array.data1[9][11] ;
 wire \data_array.data1[9][12] ;
 wire \data_array.data1[9][13] ;
 wire \data_array.data1[9][14] ;
 wire \data_array.data1[9][15] ;
 wire \data_array.data1[9][16] ;
 wire \data_array.data1[9][17] ;
 wire \data_array.data1[9][18] ;
 wire \data_array.data1[9][19] ;
 wire \data_array.data1[9][1] ;
 wire \data_array.data1[9][20] ;
 wire \data_array.data1[9][21] ;
 wire \data_array.data1[9][22] ;
 wire \data_array.data1[9][23] ;
 wire \data_array.data1[9][24] ;
 wire \data_array.data1[9][25] ;
 wire \data_array.data1[9][26] ;
 wire \data_array.data1[9][27] ;
 wire \data_array.data1[9][28] ;
 wire \data_array.data1[9][29] ;
 wire \data_array.data1[9][2] ;
 wire \data_array.data1[9][30] ;
 wire \data_array.data1[9][31] ;
 wire \data_array.data1[9][32] ;
 wire \data_array.data1[9][33] ;
 wire \data_array.data1[9][34] ;
 wire \data_array.data1[9][35] ;
 wire \data_array.data1[9][36] ;
 wire \data_array.data1[9][37] ;
 wire \data_array.data1[9][38] ;
 wire \data_array.data1[9][39] ;
 wire \data_array.data1[9][3] ;
 wire \data_array.data1[9][40] ;
 wire \data_array.data1[9][41] ;
 wire \data_array.data1[9][42] ;
 wire \data_array.data1[9][43] ;
 wire \data_array.data1[9][44] ;
 wire \data_array.data1[9][45] ;
 wire \data_array.data1[9][46] ;
 wire \data_array.data1[9][47] ;
 wire \data_array.data1[9][48] ;
 wire \data_array.data1[9][49] ;
 wire \data_array.data1[9][4] ;
 wire \data_array.data1[9][50] ;
 wire \data_array.data1[9][51] ;
 wire \data_array.data1[9][52] ;
 wire \data_array.data1[9][53] ;
 wire \data_array.data1[9][54] ;
 wire \data_array.data1[9][55] ;
 wire \data_array.data1[9][56] ;
 wire \data_array.data1[9][57] ;
 wire \data_array.data1[9][58] ;
 wire \data_array.data1[9][59] ;
 wire \data_array.data1[9][5] ;
 wire \data_array.data1[9][60] ;
 wire \data_array.data1[9][61] ;
 wire \data_array.data1[9][62] ;
 wire \data_array.data1[9][63] ;
 wire \data_array.data1[9][6] ;
 wire \data_array.data1[9][7] ;
 wire \data_array.data1[9][8] ;
 wire \data_array.data1[9][9] ;
 wire \data_array.rdata0[0] ;
 wire \data_array.rdata0[10] ;
 wire \data_array.rdata0[11] ;
 wire \data_array.rdata0[12] ;
 wire \data_array.rdata0[13] ;
 wire \data_array.rdata0[14] ;
 wire \data_array.rdata0[15] ;
 wire \data_array.rdata0[16] ;
 wire \data_array.rdata0[17] ;
 wire \data_array.rdata0[18] ;
 wire \data_array.rdata0[19] ;
 wire \data_array.rdata0[1] ;
 wire \data_array.rdata0[20] ;
 wire \data_array.rdata0[21] ;
 wire \data_array.rdata0[22] ;
 wire \data_array.rdata0[23] ;
 wire \data_array.rdata0[24] ;
 wire \data_array.rdata0[25] ;
 wire \data_array.rdata0[26] ;
 wire \data_array.rdata0[27] ;
 wire \data_array.rdata0[28] ;
 wire \data_array.rdata0[29] ;
 wire \data_array.rdata0[2] ;
 wire \data_array.rdata0[30] ;
 wire \data_array.rdata0[31] ;
 wire \data_array.rdata0[32] ;
 wire \data_array.rdata0[33] ;
 wire \data_array.rdata0[34] ;
 wire \data_array.rdata0[35] ;
 wire \data_array.rdata0[36] ;
 wire \data_array.rdata0[37] ;
 wire \data_array.rdata0[38] ;
 wire \data_array.rdata0[39] ;
 wire \data_array.rdata0[3] ;
 wire \data_array.rdata0[40] ;
 wire \data_array.rdata0[41] ;
 wire \data_array.rdata0[42] ;
 wire \data_array.rdata0[43] ;
 wire \data_array.rdata0[44] ;
 wire \data_array.rdata0[45] ;
 wire \data_array.rdata0[46] ;
 wire \data_array.rdata0[47] ;
 wire \data_array.rdata0[48] ;
 wire \data_array.rdata0[49] ;
 wire \data_array.rdata0[4] ;
 wire \data_array.rdata0[50] ;
 wire \data_array.rdata0[51] ;
 wire \data_array.rdata0[52] ;
 wire \data_array.rdata0[53] ;
 wire \data_array.rdata0[54] ;
 wire \data_array.rdata0[55] ;
 wire \data_array.rdata0[56] ;
 wire \data_array.rdata0[57] ;
 wire \data_array.rdata0[58] ;
 wire \data_array.rdata0[59] ;
 wire \data_array.rdata0[5] ;
 wire \data_array.rdata0[60] ;
 wire \data_array.rdata0[61] ;
 wire \data_array.rdata0[62] ;
 wire \data_array.rdata0[63] ;
 wire \data_array.rdata0[6] ;
 wire \data_array.rdata0[7] ;
 wire \data_array.rdata0[8] ;
 wire \data_array.rdata0[9] ;
 wire \data_array.rdata1[0] ;
 wire \data_array.rdata1[10] ;
 wire \data_array.rdata1[11] ;
 wire \data_array.rdata1[12] ;
 wire \data_array.rdata1[13] ;
 wire \data_array.rdata1[14] ;
 wire \data_array.rdata1[15] ;
 wire \data_array.rdata1[16] ;
 wire \data_array.rdata1[17] ;
 wire \data_array.rdata1[18] ;
 wire \data_array.rdata1[19] ;
 wire \data_array.rdata1[1] ;
 wire \data_array.rdata1[20] ;
 wire \data_array.rdata1[21] ;
 wire \data_array.rdata1[22] ;
 wire \data_array.rdata1[23] ;
 wire \data_array.rdata1[24] ;
 wire \data_array.rdata1[25] ;
 wire \data_array.rdata1[26] ;
 wire \data_array.rdata1[27] ;
 wire \data_array.rdata1[28] ;
 wire \data_array.rdata1[29] ;
 wire \data_array.rdata1[2] ;
 wire \data_array.rdata1[30] ;
 wire \data_array.rdata1[31] ;
 wire \data_array.rdata1[32] ;
 wire \data_array.rdata1[33] ;
 wire \data_array.rdata1[34] ;
 wire \data_array.rdata1[35] ;
 wire \data_array.rdata1[36] ;
 wire \data_array.rdata1[37] ;
 wire \data_array.rdata1[38] ;
 wire \data_array.rdata1[39] ;
 wire \data_array.rdata1[3] ;
 wire \data_array.rdata1[40] ;
 wire \data_array.rdata1[41] ;
 wire \data_array.rdata1[42] ;
 wire \data_array.rdata1[43] ;
 wire \data_array.rdata1[44] ;
 wire \data_array.rdata1[45] ;
 wire \data_array.rdata1[46] ;
 wire \data_array.rdata1[47] ;
 wire \data_array.rdata1[48] ;
 wire \data_array.rdata1[49] ;
 wire \data_array.rdata1[4] ;
 wire \data_array.rdata1[50] ;
 wire \data_array.rdata1[51] ;
 wire \data_array.rdata1[52] ;
 wire \data_array.rdata1[53] ;
 wire \data_array.rdata1[54] ;
 wire \data_array.rdata1[55] ;
 wire \data_array.rdata1[56] ;
 wire \data_array.rdata1[57] ;
 wire \data_array.rdata1[58] ;
 wire \data_array.rdata1[59] ;
 wire \data_array.rdata1[5] ;
 wire \data_array.rdata1[60] ;
 wire \data_array.rdata1[61] ;
 wire \data_array.rdata1[62] ;
 wire \data_array.rdata1[63] ;
 wire \data_array.rdata1[6] ;
 wire \data_array.rdata1[7] ;
 wire \data_array.rdata1[8] ;
 wire \data_array.rdata1[9] ;
 wire dirty_way0;
 wire dirty_way1;
 wire \fsm.lru_out ;
 wire \fsm.state[0] ;
 wire \fsm.state[2] ;
 wire \fsm.state[3] ;
 wire \fsm.state[5] ;
 wire \fsm.tag_out0[0] ;
 wire \fsm.tag_out0[10] ;
 wire \fsm.tag_out0[11] ;
 wire \fsm.tag_out0[12] ;
 wire \fsm.tag_out0[13] ;
 wire \fsm.tag_out0[14] ;
 wire \fsm.tag_out0[15] ;
 wire \fsm.tag_out0[16] ;
 wire \fsm.tag_out0[17] ;
 wire \fsm.tag_out0[18] ;
 wire \fsm.tag_out0[19] ;
 wire \fsm.tag_out0[1] ;
 wire \fsm.tag_out0[20] ;
 wire \fsm.tag_out0[21] ;
 wire \fsm.tag_out0[22] ;
 wire \fsm.tag_out0[23] ;
 wire \fsm.tag_out0[24] ;
 wire \fsm.tag_out0[2] ;
 wire \fsm.tag_out0[3] ;
 wire \fsm.tag_out0[4] ;
 wire \fsm.tag_out0[5] ;
 wire \fsm.tag_out0[6] ;
 wire \fsm.tag_out0[7] ;
 wire \fsm.tag_out0[8] ;
 wire \fsm.tag_out0[9] ;
 wire \fsm.tag_out1[0] ;
 wire \fsm.tag_out1[10] ;
 wire \fsm.tag_out1[11] ;
 wire \fsm.tag_out1[12] ;
 wire \fsm.tag_out1[13] ;
 wire \fsm.tag_out1[14] ;
 wire \fsm.tag_out1[15] ;
 wire \fsm.tag_out1[16] ;
 wire \fsm.tag_out1[17] ;
 wire \fsm.tag_out1[18] ;
 wire \fsm.tag_out1[19] ;
 wire \fsm.tag_out1[1] ;
 wire \fsm.tag_out1[20] ;
 wire \fsm.tag_out1[21] ;
 wire \fsm.tag_out1[22] ;
 wire \fsm.tag_out1[23] ;
 wire \fsm.tag_out1[24] ;
 wire \fsm.tag_out1[2] ;
 wire \fsm.tag_out1[3] ;
 wire \fsm.tag_out1[4] ;
 wire \fsm.tag_out1[5] ;
 wire \fsm.tag_out1[6] ;
 wire \fsm.tag_out1[7] ;
 wire \fsm.tag_out1[8] ;
 wire \fsm.tag_out1[9] ;
 wire \fsm.valid0 ;
 wire \fsm.valid1 ;
 wire \lru_array.lru_mem[0] ;
 wire \lru_array.lru_mem[10] ;
 wire \lru_array.lru_mem[11] ;
 wire \lru_array.lru_mem[12] ;
 wire \lru_array.lru_mem[13] ;
 wire \lru_array.lru_mem[14] ;
 wire \lru_array.lru_mem[15] ;
 wire \lru_array.lru_mem[1] ;
 wire \lru_array.lru_mem[2] ;
 wire \lru_array.lru_mem[3] ;
 wire \lru_array.lru_mem[4] ;
 wire \lru_array.lru_mem[5] ;
 wire \lru_array.lru_mem[6] ;
 wire \lru_array.lru_mem[7] ;
 wire \lru_array.lru_mem[8] ;
 wire \lru_array.lru_mem[9] ;
 wire \tag_array.dirty0[0] ;
 wire \tag_array.dirty0[10] ;
 wire \tag_array.dirty0[11] ;
 wire \tag_array.dirty0[12] ;
 wire \tag_array.dirty0[13] ;
 wire \tag_array.dirty0[14] ;
 wire \tag_array.dirty0[15] ;
 wire \tag_array.dirty0[1] ;
 wire \tag_array.dirty0[2] ;
 wire \tag_array.dirty0[3] ;
 wire \tag_array.dirty0[4] ;
 wire \tag_array.dirty0[5] ;
 wire \tag_array.dirty0[6] ;
 wire \tag_array.dirty0[7] ;
 wire \tag_array.dirty0[8] ;
 wire \tag_array.dirty0[9] ;
 wire \tag_array.dirty1[0] ;
 wire \tag_array.dirty1[10] ;
 wire \tag_array.dirty1[11] ;
 wire \tag_array.dirty1[12] ;
 wire \tag_array.dirty1[13] ;
 wire \tag_array.dirty1[14] ;
 wire \tag_array.dirty1[15] ;
 wire \tag_array.dirty1[1] ;
 wire \tag_array.dirty1[2] ;
 wire \tag_array.dirty1[3] ;
 wire \tag_array.dirty1[4] ;
 wire \tag_array.dirty1[5] ;
 wire \tag_array.dirty1[6] ;
 wire \tag_array.dirty1[7] ;
 wire \tag_array.dirty1[8] ;
 wire \tag_array.dirty1[9] ;
 wire \tag_array.tag0[0][0] ;
 wire \tag_array.tag0[0][10] ;
 wire \tag_array.tag0[0][11] ;
 wire \tag_array.tag0[0][12] ;
 wire \tag_array.tag0[0][13] ;
 wire \tag_array.tag0[0][14] ;
 wire \tag_array.tag0[0][15] ;
 wire \tag_array.tag0[0][16] ;
 wire \tag_array.tag0[0][17] ;
 wire \tag_array.tag0[0][18] ;
 wire \tag_array.tag0[0][19] ;
 wire \tag_array.tag0[0][1] ;
 wire \tag_array.tag0[0][20] ;
 wire \tag_array.tag0[0][21] ;
 wire \tag_array.tag0[0][22] ;
 wire \tag_array.tag0[0][23] ;
 wire \tag_array.tag0[0][24] ;
 wire \tag_array.tag0[0][2] ;
 wire \tag_array.tag0[0][3] ;
 wire \tag_array.tag0[0][4] ;
 wire \tag_array.tag0[0][5] ;
 wire \tag_array.tag0[0][6] ;
 wire \tag_array.tag0[0][7] ;
 wire \tag_array.tag0[0][8] ;
 wire \tag_array.tag0[0][9] ;
 wire \tag_array.tag0[10][0] ;
 wire \tag_array.tag0[10][10] ;
 wire \tag_array.tag0[10][11] ;
 wire \tag_array.tag0[10][12] ;
 wire \tag_array.tag0[10][13] ;
 wire \tag_array.tag0[10][14] ;
 wire \tag_array.tag0[10][15] ;
 wire \tag_array.tag0[10][16] ;
 wire \tag_array.tag0[10][17] ;
 wire \tag_array.tag0[10][18] ;
 wire \tag_array.tag0[10][19] ;
 wire \tag_array.tag0[10][1] ;
 wire \tag_array.tag0[10][20] ;
 wire \tag_array.tag0[10][21] ;
 wire \tag_array.tag0[10][22] ;
 wire \tag_array.tag0[10][23] ;
 wire \tag_array.tag0[10][24] ;
 wire \tag_array.tag0[10][2] ;
 wire \tag_array.tag0[10][3] ;
 wire \tag_array.tag0[10][4] ;
 wire \tag_array.tag0[10][5] ;
 wire \tag_array.tag0[10][6] ;
 wire \tag_array.tag0[10][7] ;
 wire \tag_array.tag0[10][8] ;
 wire \tag_array.tag0[10][9] ;
 wire \tag_array.tag0[11][0] ;
 wire \tag_array.tag0[11][10] ;
 wire \tag_array.tag0[11][11] ;
 wire \tag_array.tag0[11][12] ;
 wire \tag_array.tag0[11][13] ;
 wire \tag_array.tag0[11][14] ;
 wire \tag_array.tag0[11][15] ;
 wire \tag_array.tag0[11][16] ;
 wire \tag_array.tag0[11][17] ;
 wire \tag_array.tag0[11][18] ;
 wire \tag_array.tag0[11][19] ;
 wire \tag_array.tag0[11][1] ;
 wire \tag_array.tag0[11][20] ;
 wire \tag_array.tag0[11][21] ;
 wire \tag_array.tag0[11][22] ;
 wire \tag_array.tag0[11][23] ;
 wire \tag_array.tag0[11][24] ;
 wire \tag_array.tag0[11][2] ;
 wire \tag_array.tag0[11][3] ;
 wire \tag_array.tag0[11][4] ;
 wire \tag_array.tag0[11][5] ;
 wire \tag_array.tag0[11][6] ;
 wire \tag_array.tag0[11][7] ;
 wire \tag_array.tag0[11][8] ;
 wire \tag_array.tag0[11][9] ;
 wire \tag_array.tag0[12][0] ;
 wire \tag_array.tag0[12][10] ;
 wire \tag_array.tag0[12][11] ;
 wire \tag_array.tag0[12][12] ;
 wire \tag_array.tag0[12][13] ;
 wire \tag_array.tag0[12][14] ;
 wire \tag_array.tag0[12][15] ;
 wire \tag_array.tag0[12][16] ;
 wire \tag_array.tag0[12][17] ;
 wire \tag_array.tag0[12][18] ;
 wire \tag_array.tag0[12][19] ;
 wire \tag_array.tag0[12][1] ;
 wire \tag_array.tag0[12][20] ;
 wire \tag_array.tag0[12][21] ;
 wire \tag_array.tag0[12][22] ;
 wire \tag_array.tag0[12][23] ;
 wire \tag_array.tag0[12][24] ;
 wire \tag_array.tag0[12][2] ;
 wire \tag_array.tag0[12][3] ;
 wire \tag_array.tag0[12][4] ;
 wire \tag_array.tag0[12][5] ;
 wire \tag_array.tag0[12][6] ;
 wire \tag_array.tag0[12][7] ;
 wire \tag_array.tag0[12][8] ;
 wire \tag_array.tag0[12][9] ;
 wire \tag_array.tag0[13][0] ;
 wire \tag_array.tag0[13][10] ;
 wire \tag_array.tag0[13][11] ;
 wire \tag_array.tag0[13][12] ;
 wire \tag_array.tag0[13][13] ;
 wire \tag_array.tag0[13][14] ;
 wire \tag_array.tag0[13][15] ;
 wire \tag_array.tag0[13][16] ;
 wire \tag_array.tag0[13][17] ;
 wire \tag_array.tag0[13][18] ;
 wire \tag_array.tag0[13][19] ;
 wire \tag_array.tag0[13][1] ;
 wire \tag_array.tag0[13][20] ;
 wire \tag_array.tag0[13][21] ;
 wire \tag_array.tag0[13][22] ;
 wire \tag_array.tag0[13][23] ;
 wire \tag_array.tag0[13][24] ;
 wire \tag_array.tag0[13][2] ;
 wire \tag_array.tag0[13][3] ;
 wire \tag_array.tag0[13][4] ;
 wire \tag_array.tag0[13][5] ;
 wire \tag_array.tag0[13][6] ;
 wire \tag_array.tag0[13][7] ;
 wire \tag_array.tag0[13][8] ;
 wire \tag_array.tag0[13][9] ;
 wire \tag_array.tag0[14][0] ;
 wire \tag_array.tag0[14][10] ;
 wire \tag_array.tag0[14][11] ;
 wire \tag_array.tag0[14][12] ;
 wire \tag_array.tag0[14][13] ;
 wire \tag_array.tag0[14][14] ;
 wire \tag_array.tag0[14][15] ;
 wire \tag_array.tag0[14][16] ;
 wire \tag_array.tag0[14][17] ;
 wire \tag_array.tag0[14][18] ;
 wire \tag_array.tag0[14][19] ;
 wire \tag_array.tag0[14][1] ;
 wire \tag_array.tag0[14][20] ;
 wire \tag_array.tag0[14][21] ;
 wire \tag_array.tag0[14][22] ;
 wire \tag_array.tag0[14][23] ;
 wire \tag_array.tag0[14][24] ;
 wire \tag_array.tag0[14][2] ;
 wire \tag_array.tag0[14][3] ;
 wire \tag_array.tag0[14][4] ;
 wire \tag_array.tag0[14][5] ;
 wire \tag_array.tag0[14][6] ;
 wire \tag_array.tag0[14][7] ;
 wire \tag_array.tag0[14][8] ;
 wire \tag_array.tag0[14][9] ;
 wire \tag_array.tag0[15][0] ;
 wire \tag_array.tag0[15][10] ;
 wire \tag_array.tag0[15][11] ;
 wire \tag_array.tag0[15][12] ;
 wire \tag_array.tag0[15][13] ;
 wire \tag_array.tag0[15][14] ;
 wire \tag_array.tag0[15][15] ;
 wire \tag_array.tag0[15][16] ;
 wire \tag_array.tag0[15][17] ;
 wire \tag_array.tag0[15][18] ;
 wire \tag_array.tag0[15][19] ;
 wire \tag_array.tag0[15][1] ;
 wire \tag_array.tag0[15][20] ;
 wire \tag_array.tag0[15][21] ;
 wire \tag_array.tag0[15][22] ;
 wire \tag_array.tag0[15][23] ;
 wire \tag_array.tag0[15][24] ;
 wire \tag_array.tag0[15][2] ;
 wire \tag_array.tag0[15][3] ;
 wire \tag_array.tag0[15][4] ;
 wire \tag_array.tag0[15][5] ;
 wire \tag_array.tag0[15][6] ;
 wire \tag_array.tag0[15][7] ;
 wire \tag_array.tag0[15][8] ;
 wire \tag_array.tag0[15][9] ;
 wire \tag_array.tag0[1][0] ;
 wire \tag_array.tag0[1][10] ;
 wire \tag_array.tag0[1][11] ;
 wire \tag_array.tag0[1][12] ;
 wire \tag_array.tag0[1][13] ;
 wire \tag_array.tag0[1][14] ;
 wire \tag_array.tag0[1][15] ;
 wire \tag_array.tag0[1][16] ;
 wire \tag_array.tag0[1][17] ;
 wire \tag_array.tag0[1][18] ;
 wire \tag_array.tag0[1][19] ;
 wire \tag_array.tag0[1][1] ;
 wire \tag_array.tag0[1][20] ;
 wire \tag_array.tag0[1][21] ;
 wire \tag_array.tag0[1][22] ;
 wire \tag_array.tag0[1][23] ;
 wire \tag_array.tag0[1][24] ;
 wire \tag_array.tag0[1][2] ;
 wire \tag_array.tag0[1][3] ;
 wire \tag_array.tag0[1][4] ;
 wire \tag_array.tag0[1][5] ;
 wire \tag_array.tag0[1][6] ;
 wire \tag_array.tag0[1][7] ;
 wire \tag_array.tag0[1][8] ;
 wire \tag_array.tag0[1][9] ;
 wire \tag_array.tag0[2][0] ;
 wire \tag_array.tag0[2][10] ;
 wire \tag_array.tag0[2][11] ;
 wire \tag_array.tag0[2][12] ;
 wire \tag_array.tag0[2][13] ;
 wire \tag_array.tag0[2][14] ;
 wire \tag_array.tag0[2][15] ;
 wire \tag_array.tag0[2][16] ;
 wire \tag_array.tag0[2][17] ;
 wire \tag_array.tag0[2][18] ;
 wire \tag_array.tag0[2][19] ;
 wire \tag_array.tag0[2][1] ;
 wire \tag_array.tag0[2][20] ;
 wire \tag_array.tag0[2][21] ;
 wire \tag_array.tag0[2][22] ;
 wire \tag_array.tag0[2][23] ;
 wire \tag_array.tag0[2][24] ;
 wire \tag_array.tag0[2][2] ;
 wire \tag_array.tag0[2][3] ;
 wire \tag_array.tag0[2][4] ;
 wire \tag_array.tag0[2][5] ;
 wire \tag_array.tag0[2][6] ;
 wire \tag_array.tag0[2][7] ;
 wire \tag_array.tag0[2][8] ;
 wire \tag_array.tag0[2][9] ;
 wire \tag_array.tag0[3][0] ;
 wire \tag_array.tag0[3][10] ;
 wire \tag_array.tag0[3][11] ;
 wire \tag_array.tag0[3][12] ;
 wire \tag_array.tag0[3][13] ;
 wire \tag_array.tag0[3][14] ;
 wire \tag_array.tag0[3][15] ;
 wire \tag_array.tag0[3][16] ;
 wire \tag_array.tag0[3][17] ;
 wire \tag_array.tag0[3][18] ;
 wire \tag_array.tag0[3][19] ;
 wire \tag_array.tag0[3][1] ;
 wire \tag_array.tag0[3][20] ;
 wire \tag_array.tag0[3][21] ;
 wire \tag_array.tag0[3][22] ;
 wire \tag_array.tag0[3][23] ;
 wire \tag_array.tag0[3][24] ;
 wire \tag_array.tag0[3][2] ;
 wire \tag_array.tag0[3][3] ;
 wire \tag_array.tag0[3][4] ;
 wire \tag_array.tag0[3][5] ;
 wire \tag_array.tag0[3][6] ;
 wire \tag_array.tag0[3][7] ;
 wire \tag_array.tag0[3][8] ;
 wire \tag_array.tag0[3][9] ;
 wire \tag_array.tag0[4][0] ;
 wire \tag_array.tag0[4][10] ;
 wire \tag_array.tag0[4][11] ;
 wire \tag_array.tag0[4][12] ;
 wire \tag_array.tag0[4][13] ;
 wire \tag_array.tag0[4][14] ;
 wire \tag_array.tag0[4][15] ;
 wire \tag_array.tag0[4][16] ;
 wire \tag_array.tag0[4][17] ;
 wire \tag_array.tag0[4][18] ;
 wire \tag_array.tag0[4][19] ;
 wire \tag_array.tag0[4][1] ;
 wire \tag_array.tag0[4][20] ;
 wire \tag_array.tag0[4][21] ;
 wire \tag_array.tag0[4][22] ;
 wire \tag_array.tag0[4][23] ;
 wire \tag_array.tag0[4][24] ;
 wire \tag_array.tag0[4][2] ;
 wire \tag_array.tag0[4][3] ;
 wire \tag_array.tag0[4][4] ;
 wire \tag_array.tag0[4][5] ;
 wire \tag_array.tag0[4][6] ;
 wire \tag_array.tag0[4][7] ;
 wire \tag_array.tag0[4][8] ;
 wire \tag_array.tag0[4][9] ;
 wire \tag_array.tag0[5][0] ;
 wire \tag_array.tag0[5][10] ;
 wire \tag_array.tag0[5][11] ;
 wire \tag_array.tag0[5][12] ;
 wire \tag_array.tag0[5][13] ;
 wire \tag_array.tag0[5][14] ;
 wire \tag_array.tag0[5][15] ;
 wire \tag_array.tag0[5][16] ;
 wire \tag_array.tag0[5][17] ;
 wire \tag_array.tag0[5][18] ;
 wire \tag_array.tag0[5][19] ;
 wire \tag_array.tag0[5][1] ;
 wire \tag_array.tag0[5][20] ;
 wire \tag_array.tag0[5][21] ;
 wire \tag_array.tag0[5][22] ;
 wire \tag_array.tag0[5][23] ;
 wire \tag_array.tag0[5][24] ;
 wire \tag_array.tag0[5][2] ;
 wire \tag_array.tag0[5][3] ;
 wire \tag_array.tag0[5][4] ;
 wire \tag_array.tag0[5][5] ;
 wire \tag_array.tag0[5][6] ;
 wire \tag_array.tag0[5][7] ;
 wire \tag_array.tag0[5][8] ;
 wire \tag_array.tag0[5][9] ;
 wire \tag_array.tag0[6][0] ;
 wire \tag_array.tag0[6][10] ;
 wire \tag_array.tag0[6][11] ;
 wire \tag_array.tag0[6][12] ;
 wire \tag_array.tag0[6][13] ;
 wire \tag_array.tag0[6][14] ;
 wire \tag_array.tag0[6][15] ;
 wire \tag_array.tag0[6][16] ;
 wire \tag_array.tag0[6][17] ;
 wire \tag_array.tag0[6][18] ;
 wire \tag_array.tag0[6][19] ;
 wire \tag_array.tag0[6][1] ;
 wire \tag_array.tag0[6][20] ;
 wire \tag_array.tag0[6][21] ;
 wire \tag_array.tag0[6][22] ;
 wire \tag_array.tag0[6][23] ;
 wire \tag_array.tag0[6][24] ;
 wire \tag_array.tag0[6][2] ;
 wire \tag_array.tag0[6][3] ;
 wire \tag_array.tag0[6][4] ;
 wire \tag_array.tag0[6][5] ;
 wire \tag_array.tag0[6][6] ;
 wire \tag_array.tag0[6][7] ;
 wire \tag_array.tag0[6][8] ;
 wire \tag_array.tag0[6][9] ;
 wire \tag_array.tag0[7][0] ;
 wire \tag_array.tag0[7][10] ;
 wire \tag_array.tag0[7][11] ;
 wire \tag_array.tag0[7][12] ;
 wire \tag_array.tag0[7][13] ;
 wire \tag_array.tag0[7][14] ;
 wire \tag_array.tag0[7][15] ;
 wire \tag_array.tag0[7][16] ;
 wire \tag_array.tag0[7][17] ;
 wire \tag_array.tag0[7][18] ;
 wire \tag_array.tag0[7][19] ;
 wire \tag_array.tag0[7][1] ;
 wire \tag_array.tag0[7][20] ;
 wire \tag_array.tag0[7][21] ;
 wire \tag_array.tag0[7][22] ;
 wire \tag_array.tag0[7][23] ;
 wire \tag_array.tag0[7][24] ;
 wire \tag_array.tag0[7][2] ;
 wire \tag_array.tag0[7][3] ;
 wire \tag_array.tag0[7][4] ;
 wire \tag_array.tag0[7][5] ;
 wire \tag_array.tag0[7][6] ;
 wire \tag_array.tag0[7][7] ;
 wire \tag_array.tag0[7][8] ;
 wire \tag_array.tag0[7][9] ;
 wire \tag_array.tag0[8][0] ;
 wire \tag_array.tag0[8][10] ;
 wire \tag_array.tag0[8][11] ;
 wire \tag_array.tag0[8][12] ;
 wire \tag_array.tag0[8][13] ;
 wire \tag_array.tag0[8][14] ;
 wire \tag_array.tag0[8][15] ;
 wire \tag_array.tag0[8][16] ;
 wire \tag_array.tag0[8][17] ;
 wire \tag_array.tag0[8][18] ;
 wire \tag_array.tag0[8][19] ;
 wire \tag_array.tag0[8][1] ;
 wire \tag_array.tag0[8][20] ;
 wire \tag_array.tag0[8][21] ;
 wire \tag_array.tag0[8][22] ;
 wire \tag_array.tag0[8][23] ;
 wire \tag_array.tag0[8][24] ;
 wire \tag_array.tag0[8][2] ;
 wire \tag_array.tag0[8][3] ;
 wire \tag_array.tag0[8][4] ;
 wire \tag_array.tag0[8][5] ;
 wire \tag_array.tag0[8][6] ;
 wire \tag_array.tag0[8][7] ;
 wire \tag_array.tag0[8][8] ;
 wire \tag_array.tag0[8][9] ;
 wire \tag_array.tag0[9][0] ;
 wire \tag_array.tag0[9][10] ;
 wire \tag_array.tag0[9][11] ;
 wire \tag_array.tag0[9][12] ;
 wire \tag_array.tag0[9][13] ;
 wire \tag_array.tag0[9][14] ;
 wire \tag_array.tag0[9][15] ;
 wire \tag_array.tag0[9][16] ;
 wire \tag_array.tag0[9][17] ;
 wire \tag_array.tag0[9][18] ;
 wire \tag_array.tag0[9][19] ;
 wire \tag_array.tag0[9][1] ;
 wire \tag_array.tag0[9][20] ;
 wire \tag_array.tag0[9][21] ;
 wire \tag_array.tag0[9][22] ;
 wire \tag_array.tag0[9][23] ;
 wire \tag_array.tag0[9][24] ;
 wire \tag_array.tag0[9][2] ;
 wire \tag_array.tag0[9][3] ;
 wire \tag_array.tag0[9][4] ;
 wire \tag_array.tag0[9][5] ;
 wire \tag_array.tag0[9][6] ;
 wire \tag_array.tag0[9][7] ;
 wire \tag_array.tag0[9][8] ;
 wire \tag_array.tag0[9][9] ;
 wire \tag_array.tag1[0][0] ;
 wire \tag_array.tag1[0][10] ;
 wire \tag_array.tag1[0][11] ;
 wire \tag_array.tag1[0][12] ;
 wire \tag_array.tag1[0][13] ;
 wire \tag_array.tag1[0][14] ;
 wire \tag_array.tag1[0][15] ;
 wire \tag_array.tag1[0][16] ;
 wire \tag_array.tag1[0][17] ;
 wire \tag_array.tag1[0][18] ;
 wire \tag_array.tag1[0][19] ;
 wire \tag_array.tag1[0][1] ;
 wire \tag_array.tag1[0][20] ;
 wire \tag_array.tag1[0][21] ;
 wire \tag_array.tag1[0][22] ;
 wire \tag_array.tag1[0][23] ;
 wire \tag_array.tag1[0][24] ;
 wire \tag_array.tag1[0][2] ;
 wire \tag_array.tag1[0][3] ;
 wire \tag_array.tag1[0][4] ;
 wire \tag_array.tag1[0][5] ;
 wire \tag_array.tag1[0][6] ;
 wire \tag_array.tag1[0][7] ;
 wire \tag_array.tag1[0][8] ;
 wire \tag_array.tag1[0][9] ;
 wire \tag_array.tag1[10][0] ;
 wire \tag_array.tag1[10][10] ;
 wire \tag_array.tag1[10][11] ;
 wire \tag_array.tag1[10][12] ;
 wire \tag_array.tag1[10][13] ;
 wire \tag_array.tag1[10][14] ;
 wire \tag_array.tag1[10][15] ;
 wire \tag_array.tag1[10][16] ;
 wire \tag_array.tag1[10][17] ;
 wire \tag_array.tag1[10][18] ;
 wire \tag_array.tag1[10][19] ;
 wire \tag_array.tag1[10][1] ;
 wire \tag_array.tag1[10][20] ;
 wire \tag_array.tag1[10][21] ;
 wire \tag_array.tag1[10][22] ;
 wire \tag_array.tag1[10][23] ;
 wire \tag_array.tag1[10][24] ;
 wire \tag_array.tag1[10][2] ;
 wire \tag_array.tag1[10][3] ;
 wire \tag_array.tag1[10][4] ;
 wire \tag_array.tag1[10][5] ;
 wire \tag_array.tag1[10][6] ;
 wire \tag_array.tag1[10][7] ;
 wire \tag_array.tag1[10][8] ;
 wire \tag_array.tag1[10][9] ;
 wire \tag_array.tag1[11][0] ;
 wire \tag_array.tag1[11][10] ;
 wire \tag_array.tag1[11][11] ;
 wire \tag_array.tag1[11][12] ;
 wire \tag_array.tag1[11][13] ;
 wire \tag_array.tag1[11][14] ;
 wire \tag_array.tag1[11][15] ;
 wire \tag_array.tag1[11][16] ;
 wire \tag_array.tag1[11][17] ;
 wire \tag_array.tag1[11][18] ;
 wire \tag_array.tag1[11][19] ;
 wire \tag_array.tag1[11][1] ;
 wire \tag_array.tag1[11][20] ;
 wire \tag_array.tag1[11][21] ;
 wire \tag_array.tag1[11][22] ;
 wire \tag_array.tag1[11][23] ;
 wire \tag_array.tag1[11][24] ;
 wire \tag_array.tag1[11][2] ;
 wire \tag_array.tag1[11][3] ;
 wire \tag_array.tag1[11][4] ;
 wire \tag_array.tag1[11][5] ;
 wire \tag_array.tag1[11][6] ;
 wire \tag_array.tag1[11][7] ;
 wire \tag_array.tag1[11][8] ;
 wire \tag_array.tag1[11][9] ;
 wire \tag_array.tag1[12][0] ;
 wire \tag_array.tag1[12][10] ;
 wire \tag_array.tag1[12][11] ;
 wire \tag_array.tag1[12][12] ;
 wire \tag_array.tag1[12][13] ;
 wire \tag_array.tag1[12][14] ;
 wire \tag_array.tag1[12][15] ;
 wire \tag_array.tag1[12][16] ;
 wire \tag_array.tag1[12][17] ;
 wire \tag_array.tag1[12][18] ;
 wire \tag_array.tag1[12][19] ;
 wire \tag_array.tag1[12][1] ;
 wire \tag_array.tag1[12][20] ;
 wire \tag_array.tag1[12][21] ;
 wire \tag_array.tag1[12][22] ;
 wire \tag_array.tag1[12][23] ;
 wire \tag_array.tag1[12][24] ;
 wire \tag_array.tag1[12][2] ;
 wire \tag_array.tag1[12][3] ;
 wire \tag_array.tag1[12][4] ;
 wire \tag_array.tag1[12][5] ;
 wire \tag_array.tag1[12][6] ;
 wire \tag_array.tag1[12][7] ;
 wire \tag_array.tag1[12][8] ;
 wire \tag_array.tag1[12][9] ;
 wire \tag_array.tag1[13][0] ;
 wire \tag_array.tag1[13][10] ;
 wire \tag_array.tag1[13][11] ;
 wire \tag_array.tag1[13][12] ;
 wire \tag_array.tag1[13][13] ;
 wire \tag_array.tag1[13][14] ;
 wire \tag_array.tag1[13][15] ;
 wire \tag_array.tag1[13][16] ;
 wire \tag_array.tag1[13][17] ;
 wire \tag_array.tag1[13][18] ;
 wire \tag_array.tag1[13][19] ;
 wire \tag_array.tag1[13][1] ;
 wire \tag_array.tag1[13][20] ;
 wire \tag_array.tag1[13][21] ;
 wire \tag_array.tag1[13][22] ;
 wire \tag_array.tag1[13][23] ;
 wire \tag_array.tag1[13][24] ;
 wire \tag_array.tag1[13][2] ;
 wire \tag_array.tag1[13][3] ;
 wire \tag_array.tag1[13][4] ;
 wire \tag_array.tag1[13][5] ;
 wire \tag_array.tag1[13][6] ;
 wire \tag_array.tag1[13][7] ;
 wire \tag_array.tag1[13][8] ;
 wire \tag_array.tag1[13][9] ;
 wire \tag_array.tag1[14][0] ;
 wire \tag_array.tag1[14][10] ;
 wire \tag_array.tag1[14][11] ;
 wire \tag_array.tag1[14][12] ;
 wire \tag_array.tag1[14][13] ;
 wire \tag_array.tag1[14][14] ;
 wire \tag_array.tag1[14][15] ;
 wire \tag_array.tag1[14][16] ;
 wire \tag_array.tag1[14][17] ;
 wire \tag_array.tag1[14][18] ;
 wire \tag_array.tag1[14][19] ;
 wire \tag_array.tag1[14][1] ;
 wire \tag_array.tag1[14][20] ;
 wire \tag_array.tag1[14][21] ;
 wire \tag_array.tag1[14][22] ;
 wire \tag_array.tag1[14][23] ;
 wire \tag_array.tag1[14][24] ;
 wire \tag_array.tag1[14][2] ;
 wire \tag_array.tag1[14][3] ;
 wire \tag_array.tag1[14][4] ;
 wire \tag_array.tag1[14][5] ;
 wire \tag_array.tag1[14][6] ;
 wire \tag_array.tag1[14][7] ;
 wire \tag_array.tag1[14][8] ;
 wire \tag_array.tag1[14][9] ;
 wire \tag_array.tag1[15][0] ;
 wire \tag_array.tag1[15][10] ;
 wire \tag_array.tag1[15][11] ;
 wire \tag_array.tag1[15][12] ;
 wire \tag_array.tag1[15][13] ;
 wire \tag_array.tag1[15][14] ;
 wire \tag_array.tag1[15][15] ;
 wire \tag_array.tag1[15][16] ;
 wire \tag_array.tag1[15][17] ;
 wire \tag_array.tag1[15][18] ;
 wire \tag_array.tag1[15][19] ;
 wire \tag_array.tag1[15][1] ;
 wire \tag_array.tag1[15][20] ;
 wire \tag_array.tag1[15][21] ;
 wire \tag_array.tag1[15][22] ;
 wire \tag_array.tag1[15][23] ;
 wire \tag_array.tag1[15][24] ;
 wire \tag_array.tag1[15][2] ;
 wire \tag_array.tag1[15][3] ;
 wire \tag_array.tag1[15][4] ;
 wire \tag_array.tag1[15][5] ;
 wire \tag_array.tag1[15][6] ;
 wire \tag_array.tag1[15][7] ;
 wire \tag_array.tag1[15][8] ;
 wire \tag_array.tag1[15][9] ;
 wire \tag_array.tag1[1][0] ;
 wire \tag_array.tag1[1][10] ;
 wire \tag_array.tag1[1][11] ;
 wire \tag_array.tag1[1][12] ;
 wire \tag_array.tag1[1][13] ;
 wire \tag_array.tag1[1][14] ;
 wire \tag_array.tag1[1][15] ;
 wire \tag_array.tag1[1][16] ;
 wire \tag_array.tag1[1][17] ;
 wire \tag_array.tag1[1][18] ;
 wire \tag_array.tag1[1][19] ;
 wire \tag_array.tag1[1][1] ;
 wire \tag_array.tag1[1][20] ;
 wire \tag_array.tag1[1][21] ;
 wire \tag_array.tag1[1][22] ;
 wire \tag_array.tag1[1][23] ;
 wire \tag_array.tag1[1][24] ;
 wire \tag_array.tag1[1][2] ;
 wire \tag_array.tag1[1][3] ;
 wire \tag_array.tag1[1][4] ;
 wire \tag_array.tag1[1][5] ;
 wire \tag_array.tag1[1][6] ;
 wire \tag_array.tag1[1][7] ;
 wire \tag_array.tag1[1][8] ;
 wire \tag_array.tag1[1][9] ;
 wire \tag_array.tag1[2][0] ;
 wire \tag_array.tag1[2][10] ;
 wire \tag_array.tag1[2][11] ;
 wire \tag_array.tag1[2][12] ;
 wire \tag_array.tag1[2][13] ;
 wire \tag_array.tag1[2][14] ;
 wire \tag_array.tag1[2][15] ;
 wire \tag_array.tag1[2][16] ;
 wire \tag_array.tag1[2][17] ;
 wire \tag_array.tag1[2][18] ;
 wire \tag_array.tag1[2][19] ;
 wire \tag_array.tag1[2][1] ;
 wire \tag_array.tag1[2][20] ;
 wire \tag_array.tag1[2][21] ;
 wire \tag_array.tag1[2][22] ;
 wire \tag_array.tag1[2][23] ;
 wire \tag_array.tag1[2][24] ;
 wire \tag_array.tag1[2][2] ;
 wire \tag_array.tag1[2][3] ;
 wire \tag_array.tag1[2][4] ;
 wire \tag_array.tag1[2][5] ;
 wire \tag_array.tag1[2][6] ;
 wire \tag_array.tag1[2][7] ;
 wire \tag_array.tag1[2][8] ;
 wire \tag_array.tag1[2][9] ;
 wire \tag_array.tag1[3][0] ;
 wire \tag_array.tag1[3][10] ;
 wire \tag_array.tag1[3][11] ;
 wire \tag_array.tag1[3][12] ;
 wire \tag_array.tag1[3][13] ;
 wire \tag_array.tag1[3][14] ;
 wire \tag_array.tag1[3][15] ;
 wire \tag_array.tag1[3][16] ;
 wire \tag_array.tag1[3][17] ;
 wire \tag_array.tag1[3][18] ;
 wire \tag_array.tag1[3][19] ;
 wire \tag_array.tag1[3][1] ;
 wire \tag_array.tag1[3][20] ;
 wire \tag_array.tag1[3][21] ;
 wire \tag_array.tag1[3][22] ;
 wire \tag_array.tag1[3][23] ;
 wire \tag_array.tag1[3][24] ;
 wire \tag_array.tag1[3][2] ;
 wire \tag_array.tag1[3][3] ;
 wire \tag_array.tag1[3][4] ;
 wire \tag_array.tag1[3][5] ;
 wire \tag_array.tag1[3][6] ;
 wire \tag_array.tag1[3][7] ;
 wire \tag_array.tag1[3][8] ;
 wire \tag_array.tag1[3][9] ;
 wire \tag_array.tag1[4][0] ;
 wire \tag_array.tag1[4][10] ;
 wire \tag_array.tag1[4][11] ;
 wire \tag_array.tag1[4][12] ;
 wire \tag_array.tag1[4][13] ;
 wire \tag_array.tag1[4][14] ;
 wire \tag_array.tag1[4][15] ;
 wire \tag_array.tag1[4][16] ;
 wire \tag_array.tag1[4][17] ;
 wire \tag_array.tag1[4][18] ;
 wire \tag_array.tag1[4][19] ;
 wire \tag_array.tag1[4][1] ;
 wire \tag_array.tag1[4][20] ;
 wire \tag_array.tag1[4][21] ;
 wire \tag_array.tag1[4][22] ;
 wire \tag_array.tag1[4][23] ;
 wire \tag_array.tag1[4][24] ;
 wire \tag_array.tag1[4][2] ;
 wire \tag_array.tag1[4][3] ;
 wire \tag_array.tag1[4][4] ;
 wire \tag_array.tag1[4][5] ;
 wire \tag_array.tag1[4][6] ;
 wire \tag_array.tag1[4][7] ;
 wire \tag_array.tag1[4][8] ;
 wire \tag_array.tag1[4][9] ;
 wire \tag_array.tag1[5][0] ;
 wire \tag_array.tag1[5][10] ;
 wire \tag_array.tag1[5][11] ;
 wire \tag_array.tag1[5][12] ;
 wire \tag_array.tag1[5][13] ;
 wire \tag_array.tag1[5][14] ;
 wire \tag_array.tag1[5][15] ;
 wire \tag_array.tag1[5][16] ;
 wire \tag_array.tag1[5][17] ;
 wire \tag_array.tag1[5][18] ;
 wire \tag_array.tag1[5][19] ;
 wire \tag_array.tag1[5][1] ;
 wire \tag_array.tag1[5][20] ;
 wire \tag_array.tag1[5][21] ;
 wire \tag_array.tag1[5][22] ;
 wire \tag_array.tag1[5][23] ;
 wire \tag_array.tag1[5][24] ;
 wire \tag_array.tag1[5][2] ;
 wire \tag_array.tag1[5][3] ;
 wire \tag_array.tag1[5][4] ;
 wire \tag_array.tag1[5][5] ;
 wire \tag_array.tag1[5][6] ;
 wire \tag_array.tag1[5][7] ;
 wire \tag_array.tag1[5][8] ;
 wire \tag_array.tag1[5][9] ;
 wire \tag_array.tag1[6][0] ;
 wire \tag_array.tag1[6][10] ;
 wire \tag_array.tag1[6][11] ;
 wire \tag_array.tag1[6][12] ;
 wire \tag_array.tag1[6][13] ;
 wire \tag_array.tag1[6][14] ;
 wire \tag_array.tag1[6][15] ;
 wire \tag_array.tag1[6][16] ;
 wire \tag_array.tag1[6][17] ;
 wire \tag_array.tag1[6][18] ;
 wire \tag_array.tag1[6][19] ;
 wire \tag_array.tag1[6][1] ;
 wire \tag_array.tag1[6][20] ;
 wire \tag_array.tag1[6][21] ;
 wire \tag_array.tag1[6][22] ;
 wire \tag_array.tag1[6][23] ;
 wire \tag_array.tag1[6][24] ;
 wire \tag_array.tag1[6][2] ;
 wire \tag_array.tag1[6][3] ;
 wire \tag_array.tag1[6][4] ;
 wire \tag_array.tag1[6][5] ;
 wire \tag_array.tag1[6][6] ;
 wire \tag_array.tag1[6][7] ;
 wire \tag_array.tag1[6][8] ;
 wire \tag_array.tag1[6][9] ;
 wire \tag_array.tag1[7][0] ;
 wire \tag_array.tag1[7][10] ;
 wire \tag_array.tag1[7][11] ;
 wire \tag_array.tag1[7][12] ;
 wire \tag_array.tag1[7][13] ;
 wire \tag_array.tag1[7][14] ;
 wire \tag_array.tag1[7][15] ;
 wire \tag_array.tag1[7][16] ;
 wire \tag_array.tag1[7][17] ;
 wire \tag_array.tag1[7][18] ;
 wire \tag_array.tag1[7][19] ;
 wire \tag_array.tag1[7][1] ;
 wire \tag_array.tag1[7][20] ;
 wire \tag_array.tag1[7][21] ;
 wire \tag_array.tag1[7][22] ;
 wire \tag_array.tag1[7][23] ;
 wire \tag_array.tag1[7][24] ;
 wire \tag_array.tag1[7][2] ;
 wire \tag_array.tag1[7][3] ;
 wire \tag_array.tag1[7][4] ;
 wire \tag_array.tag1[7][5] ;
 wire \tag_array.tag1[7][6] ;
 wire \tag_array.tag1[7][7] ;
 wire \tag_array.tag1[7][8] ;
 wire \tag_array.tag1[7][9] ;
 wire \tag_array.tag1[8][0] ;
 wire \tag_array.tag1[8][10] ;
 wire \tag_array.tag1[8][11] ;
 wire \tag_array.tag1[8][12] ;
 wire \tag_array.tag1[8][13] ;
 wire \tag_array.tag1[8][14] ;
 wire \tag_array.tag1[8][15] ;
 wire \tag_array.tag1[8][16] ;
 wire \tag_array.tag1[8][17] ;
 wire \tag_array.tag1[8][18] ;
 wire \tag_array.tag1[8][19] ;
 wire \tag_array.tag1[8][1] ;
 wire \tag_array.tag1[8][20] ;
 wire \tag_array.tag1[8][21] ;
 wire \tag_array.tag1[8][22] ;
 wire \tag_array.tag1[8][23] ;
 wire \tag_array.tag1[8][24] ;
 wire \tag_array.tag1[8][2] ;
 wire \tag_array.tag1[8][3] ;
 wire \tag_array.tag1[8][4] ;
 wire \tag_array.tag1[8][5] ;
 wire \tag_array.tag1[8][6] ;
 wire \tag_array.tag1[8][7] ;
 wire \tag_array.tag1[8][8] ;
 wire \tag_array.tag1[8][9] ;
 wire \tag_array.tag1[9][0] ;
 wire \tag_array.tag1[9][10] ;
 wire \tag_array.tag1[9][11] ;
 wire \tag_array.tag1[9][12] ;
 wire \tag_array.tag1[9][13] ;
 wire \tag_array.tag1[9][14] ;
 wire \tag_array.tag1[9][15] ;
 wire \tag_array.tag1[9][16] ;
 wire \tag_array.tag1[9][17] ;
 wire \tag_array.tag1[9][18] ;
 wire \tag_array.tag1[9][19] ;
 wire \tag_array.tag1[9][1] ;
 wire \tag_array.tag1[9][20] ;
 wire \tag_array.tag1[9][21] ;
 wire \tag_array.tag1[9][22] ;
 wire \tag_array.tag1[9][23] ;
 wire \tag_array.tag1[9][24] ;
 wire \tag_array.tag1[9][2] ;
 wire \tag_array.tag1[9][3] ;
 wire \tag_array.tag1[9][4] ;
 wire \tag_array.tag1[9][5] ;
 wire \tag_array.tag1[9][6] ;
 wire \tag_array.tag1[9][7] ;
 wire \tag_array.tag1[9][8] ;
 wire \tag_array.tag1[9][9] ;
 wire \tag_array.valid0[0] ;
 wire \tag_array.valid0[10] ;
 wire \tag_array.valid0[11] ;
 wire \tag_array.valid0[12] ;
 wire \tag_array.valid0[13] ;
 wire \tag_array.valid0[14] ;
 wire \tag_array.valid0[15] ;
 wire \tag_array.valid0[1] ;
 wire \tag_array.valid0[2] ;
 wire \tag_array.valid0[3] ;
 wire \tag_array.valid0[4] ;
 wire \tag_array.valid0[5] ;
 wire \tag_array.valid0[6] ;
 wire \tag_array.valid0[7] ;
 wire \tag_array.valid0[8] ;
 wire \tag_array.valid0[9] ;
 wire \tag_array.valid1[0] ;
 wire \tag_array.valid1[10] ;
 wire \tag_array.valid1[11] ;
 wire \tag_array.valid1[12] ;
 wire \tag_array.valid1[13] ;
 wire \tag_array.valid1[14] ;
 wire \tag_array.valid1[15] ;
 wire \tag_array.valid1[1] ;
 wire \tag_array.valid1[2] ;
 wire \tag_array.valid1[3] ;
 wire \tag_array.valid1[4] ;
 wire \tag_array.valid1[5] ;
 wire \tag_array.valid1[6] ;
 wire \tag_array.valid1[7] ;
 wire \tag_array.valid1[8] ;
 wire \tag_array.valid1[9] ;

 sky130_fd_sc_hd__inv_2 _05612_ (.A(mem_ready),
    .Y(_03134_));
 sky130_fd_sc_hd__inv_2 _05613_ (.A(cpu_addr[8]),
    .Y(_03135_));
 sky130_fd_sc_hd__inv_2 _05614_ (.A(cpu_addr[9]),
    .Y(_03136_));
 sky130_fd_sc_hd__inv_2 _05615_ (.A(\fsm.tag_out1[3] ),
    .Y(_03137_));
 sky130_fd_sc_hd__inv_2 _05616_ (.A(\fsm.tag_out1[6] ),
    .Y(_03138_));
 sky130_fd_sc_hd__inv_2 _05617_ (.A(cpu_addr[18]),
    .Y(_03139_));
 sky130_fd_sc_hd__inv_2 _05618_ (.A(cpu_addr[21]),
    .Y(_03140_));
 sky130_fd_sc_hd__inv_2 _05619_ (.A(\fsm.tag_out1[15] ),
    .Y(_03141_));
 sky130_fd_sc_hd__inv_2 _05620_ (.A(cpu_addr[25]),
    .Y(_03142_));
 sky130_fd_sc_hd__inv_2 _05621_ (.A(cpu_addr[27]),
    .Y(_03143_));
 sky130_fd_sc_hd__inv_2 _05622_ (.A(\fsm.tag_out1[20] ),
    .Y(_03144_));
 sky130_fd_sc_hd__inv_2 _05623_ (.A(\fsm.tag_out0[18] ),
    .Y(_03145_));
 sky130_fd_sc_hd__inv_2 _05624_ (.A(reset),
    .Y(_00189_));
 sky130_fd_sc_hd__and2_2 _05625_ (.A(mem_ready),
    .B(mem_read),
    .X(_03146_));
 sky130_fd_sc_hd__nand2_2 _05626_ (.A(mem_ready),
    .B(mem_read),
    .Y(_03147_));
 sky130_fd_sc_hd__or2_2 _05627_ (.A(\fsm.state[2] ),
    .B(_03146_),
    .X(cpu_ready));
 sky130_fd_sc_hd__nor2_2 _05628_ (.A(cpu_write),
    .B(cpu_read),
    .Y(_03148_));
 sky130_fd_sc_hd__a21o_2 _05629_ (.A1(\fsm.state[0] ),
    .A2(_03148_),
    .B1(cpu_ready),
    .X(_00186_));
 sky130_fd_sc_hd__and3b_2 _05630_ (.A_N(\fsm.lru_out ),
    .B(dirty_way0),
    .C(\fsm.valid0 ),
    .X(_03149_));
 sky130_fd_sc_hd__a31o_2 _05631_ (.A1(\fsm.lru_out ),
    .A2(\fsm.valid1 ),
    .A3(dirty_way1),
    .B1(_03149_),
    .X(_03150_));
 sky130_fd_sc_hd__inv_2 _05632_ (.A(_03150_),
    .Y(_03151_));
 sky130_fd_sc_hd__mux2_1 _05633_ (.A0(mem_read),
    .A1(mem_write),
    .S(mem_ready),
    .X(_03152_));
 sky130_fd_sc_hd__a21o_2 _05634_ (.A1(\fsm.state[5] ),
    .A2(_03151_),
    .B1(_03152_),
    .X(_00188_));
 sky130_fd_sc_hd__a22o_2 _05635_ (.A1(_03134_),
    .A2(mem_write),
    .B1(_03150_),
    .B2(\fsm.state[5] ),
    .X(_00187_));
 sky130_fd_sc_hd__and3_2 _05636_ (.A(mem_ready),
    .B(mem_read),
    .C(cpu_read),
    .X(_03153_));
 sky130_fd_sc_hd__and2_2 _05637_ (.A(\fsm.state[2] ),
    .B(cpu_read),
    .X(_03154_));
 sky130_fd_sc_hd__xor2_2 _05638_ (.A(cpu_addr[19]),
    .B(\fsm.tag_out0[12] ),
    .X(_03155_));
 sky130_fd_sc_hd__xor2_2 _05639_ (.A(cpu_addr[31]),
    .B(\fsm.tag_out0[24] ),
    .X(_03156_));
 sky130_fd_sc_hd__xor2_2 _05640_ (.A(cpu_addr[25]),
    .B(\fsm.tag_out0[18] ),
    .X(_03157_));
 sky130_fd_sc_hd__xor2_2 _05641_ (.A(cpu_addr[15]),
    .B(\fsm.tag_out0[8] ),
    .X(_03158_));
 sky130_fd_sc_hd__or4_2 _05642_ (.A(_03155_),
    .B(_03156_),
    .C(_03157_),
    .D(_03158_),
    .X(_03159_));
 sky130_fd_sc_hd__and2b_2 _05643_ (.A_N(cpu_addr[7]),
    .B(\fsm.tag_out0[0] ),
    .X(_03160_));
 sky130_fd_sc_hd__xor2_2 _05644_ (.A(cpu_addr[8]),
    .B(\fsm.tag_out0[1] ),
    .X(_03161_));
 sky130_fd_sc_hd__or3b_2 _05645_ (.A(_03160_),
    .B(_03161_),
    .C_N(\fsm.valid0 ),
    .X(_03162_));
 sky130_fd_sc_hd__xor2_2 _05646_ (.A(cpu_addr[30]),
    .B(\fsm.tag_out0[23] ),
    .X(_03163_));
 sky130_fd_sc_hd__nand2_2 _05647_ (.A(cpu_addr[9]),
    .B(\fsm.tag_out0[2] ),
    .Y(_03164_));
 sky130_fd_sc_hd__or2_2 _05648_ (.A(cpu_addr[9]),
    .B(\fsm.tag_out0[2] ),
    .X(_03165_));
 sky130_fd_sc_hd__a21o_2 _05649_ (.A1(_03164_),
    .A2(_03165_),
    .B1(_03163_),
    .X(_03166_));
 sky130_fd_sc_hd__and2b_2 _05650_ (.A_N(cpu_addr[27]),
    .B(\fsm.tag_out0[20] ),
    .X(_03167_));
 sky130_fd_sc_hd__and2b_2 _05651_ (.A_N(\fsm.tag_out0[0] ),
    .B(cpu_addr[7]),
    .X(_03168_));
 sky130_fd_sc_hd__and2b_2 _05652_ (.A_N(cpu_addr[11]),
    .B(\fsm.tag_out0[4] ),
    .X(_03169_));
 sky130_fd_sc_hd__and2b_2 _05653_ (.A_N(\fsm.tag_out0[3] ),
    .B(cpu_addr[10]),
    .X(_03170_));
 sky130_fd_sc_hd__or4_2 _05654_ (.A(_03167_),
    .B(_03168_),
    .C(_03169_),
    .D(_03170_),
    .X(_03171_));
 sky130_fd_sc_hd__and2b_2 _05655_ (.A_N(\fsm.tag_out0[21] ),
    .B(cpu_addr[28]),
    .X(_03172_));
 sky130_fd_sc_hd__and2b_2 _05656_ (.A_N(\fsm.tag_out0[11] ),
    .B(cpu_addr[18]),
    .X(_03173_));
 sky130_fd_sc_hd__and2b_2 _05657_ (.A_N(cpu_addr[12]),
    .B(\fsm.tag_out0[5] ),
    .X(_03174_));
 sky130_fd_sc_hd__and2b_2 _05658_ (.A_N(\fsm.tag_out0[19] ),
    .B(cpu_addr[26]),
    .X(_03175_));
 sky130_fd_sc_hd__or4_2 _05659_ (.A(_03172_),
    .B(_03173_),
    .C(_03174_),
    .D(_03175_),
    .X(_03176_));
 sky130_fd_sc_hd__or4_2 _05660_ (.A(_03162_),
    .B(_03166_),
    .C(_03171_),
    .D(_03176_),
    .X(_03177_));
 sky130_fd_sc_hd__and2b_2 _05661_ (.A_N(cpu_addr[23]),
    .B(\fsm.tag_out0[16] ),
    .X(_03178_));
 sky130_fd_sc_hd__and2b_2 _05662_ (.A_N(cpu_addr[22]),
    .B(\fsm.tag_out0[15] ),
    .X(_03179_));
 sky130_fd_sc_hd__and2b_2 _05663_ (.A_N(cpu_addr[10]),
    .B(\fsm.tag_out0[3] ),
    .X(_03180_));
 sky130_fd_sc_hd__or3_2 _05664_ (.A(_03178_),
    .B(_03179_),
    .C(_03180_),
    .X(_03181_));
 sky130_fd_sc_hd__and2b_2 _05665_ (.A_N(\fsm.tag_out0[4] ),
    .B(cpu_addr[11]),
    .X(_03182_));
 sky130_fd_sc_hd__and2b_2 _05666_ (.A_N(cpu_addr[14]),
    .B(\fsm.tag_out0[7] ),
    .X(_03183_));
 sky130_fd_sc_hd__and2b_2 _05667_ (.A_N(\fsm.tag_out0[16] ),
    .B(cpu_addr[23]),
    .X(_03184_));
 sky130_fd_sc_hd__and2b_2 _05668_ (.A_N(cpu_addr[18]),
    .B(\fsm.tag_out0[11] ),
    .X(_03185_));
 sky130_fd_sc_hd__or4_2 _05669_ (.A(_03182_),
    .B(_03183_),
    .C(_03184_),
    .D(_03185_),
    .X(_03186_));
 sky130_fd_sc_hd__and2b_2 _05670_ (.A_N(\fsm.tag_out0[10] ),
    .B(cpu_addr[17]),
    .X(_03187_));
 sky130_fd_sc_hd__and2b_2 _05671_ (.A_N(cpu_addr[21]),
    .B(\fsm.tag_out0[14] ),
    .X(_03188_));
 sky130_fd_sc_hd__and2b_2 _05672_ (.A_N(\fsm.tag_out0[15] ),
    .B(cpu_addr[22]),
    .X(_03189_));
 sky130_fd_sc_hd__and2b_2 _05673_ (.A_N(\fsm.tag_out0[14] ),
    .B(cpu_addr[21]),
    .X(_03190_));
 sky130_fd_sc_hd__or4_2 _05674_ (.A(_03187_),
    .B(_03188_),
    .C(_03189_),
    .D(_03190_),
    .X(_03191_));
 sky130_fd_sc_hd__or3_2 _05675_ (.A(_03181_),
    .B(_03186_),
    .C(_03191_),
    .X(_03192_));
 sky130_fd_sc_hd__and2b_2 _05676_ (.A_N(\fsm.tag_out0[20] ),
    .B(cpu_addr[27]),
    .X(_03193_));
 sky130_fd_sc_hd__and2b_2 _05677_ (.A_N(\fsm.tag_out0[9] ),
    .B(cpu_addr[16]),
    .X(_03194_));
 sky130_fd_sc_hd__and2b_2 _05678_ (.A_N(cpu_addr[13]),
    .B(\fsm.tag_out0[6] ),
    .X(_03195_));
 sky130_fd_sc_hd__and2b_2 _05679_ (.A_N(\fsm.tag_out0[6] ),
    .B(cpu_addr[13]),
    .X(_03196_));
 sky130_fd_sc_hd__or4_2 _05680_ (.A(_03193_),
    .B(_03194_),
    .C(_03195_),
    .D(_03196_),
    .X(_03197_));
 sky130_fd_sc_hd__and2b_2 _05681_ (.A_N(cpu_addr[17]),
    .B(\fsm.tag_out0[10] ),
    .X(_03198_));
 sky130_fd_sc_hd__and2b_2 _05682_ (.A_N(\fsm.tag_out0[5] ),
    .B(cpu_addr[12]),
    .X(_03199_));
 sky130_fd_sc_hd__and2b_2 _05683_ (.A_N(cpu_addr[29]),
    .B(\fsm.tag_out0[22] ),
    .X(_03200_));
 sky130_fd_sc_hd__and2b_2 _05684_ (.A_N(cpu_addr[16]),
    .B(\fsm.tag_out0[9] ),
    .X(_03201_));
 sky130_fd_sc_hd__or4_2 _05685_ (.A(_03198_),
    .B(_03199_),
    .C(_03200_),
    .D(_03201_),
    .X(_03202_));
 sky130_fd_sc_hd__xor2_2 _05686_ (.A(cpu_addr[20]),
    .B(\fsm.tag_out0[13] ),
    .X(_03203_));
 sky130_fd_sc_hd__and2b_2 _05687_ (.A_N(cpu_addr[24]),
    .B(\fsm.tag_out0[17] ),
    .X(_03204_));
 sky130_fd_sc_hd__and2b_2 _05688_ (.A_N(\fsm.tag_out0[17] ),
    .B(cpu_addr[24]),
    .X(_03205_));
 sky130_fd_sc_hd__or3_2 _05689_ (.A(_03203_),
    .B(_03204_),
    .C(_03205_),
    .X(_03206_));
 sky130_fd_sc_hd__and2b_2 _05690_ (.A_N(cpu_addr[26]),
    .B(\fsm.tag_out0[19] ),
    .X(_03207_));
 sky130_fd_sc_hd__and2b_2 _05691_ (.A_N(\fsm.tag_out0[7] ),
    .B(cpu_addr[14]),
    .X(_03208_));
 sky130_fd_sc_hd__and2b_2 _05692_ (.A_N(\fsm.tag_out0[22] ),
    .B(cpu_addr[29]),
    .X(_03209_));
 sky130_fd_sc_hd__and2b_2 _05693_ (.A_N(cpu_addr[28]),
    .B(\fsm.tag_out0[21] ),
    .X(_03210_));
 sky130_fd_sc_hd__or4_2 _05694_ (.A(_03207_),
    .B(_03208_),
    .C(_03209_),
    .D(_03210_),
    .X(_03211_));
 sky130_fd_sc_hd__or4_2 _05695_ (.A(_03197_),
    .B(_03202_),
    .C(_03206_),
    .D(_03211_),
    .X(_03212_));
 sky130_fd_sc_hd__or4_2 _05696_ (.A(_03159_),
    .B(_03177_),
    .C(_03192_),
    .D(_03212_),
    .X(_03213_));
 sky130_fd_sc_hd__or2_2 _05697_ (.A(_03167_),
    .B(_03193_),
    .X(_03214_));
 sky130_fd_sc_hd__a211o_2 _05698_ (.A1(cpu_addr[25]),
    .A2(_03145_),
    .B1(_03155_),
    .C1(_03209_),
    .X(_03215_));
 sky130_fd_sc_hd__a2111o_2 _05699_ (.A1(_03142_),
    .A2(\fsm.tag_out0[18] ),
    .B1(_03172_),
    .C1(_03178_),
    .D1(_03207_),
    .X(_03216_));
 sky130_fd_sc_hd__or3_2 _05700_ (.A(_03214_),
    .B(_03215_),
    .C(_03216_),
    .X(_03217_));
 sky130_fd_sc_hd__and2b_2 _05701_ (.A_N(\fsm.tag_out0[1] ),
    .B(cpu_addr[8]),
    .X(_03218_));
 sky130_fd_sc_hd__or3_2 _05702_ (.A(_03187_),
    .B(_03188_),
    .C(_03218_),
    .X(_03219_));
 sky130_fd_sc_hd__nand2_2 _05703_ (.A(cpu_addr[7]),
    .B(\fsm.tag_out0[0] ),
    .Y(_03220_));
 sky130_fd_sc_hd__or2_2 _05704_ (.A(cpu_addr[7]),
    .B(\fsm.tag_out0[0] ),
    .X(_03221_));
 sky130_fd_sc_hd__a211o_2 _05705_ (.A1(_03220_),
    .A2(_03221_),
    .B1(_03180_),
    .C1(_03210_),
    .X(_03222_));
 sky130_fd_sc_hd__or3_2 _05706_ (.A(_03163_),
    .B(_03183_),
    .C(_03201_),
    .X(_03223_));
 sky130_fd_sc_hd__and2b_2 _05707_ (.A_N(cpu_addr[9]),
    .B(\fsm.tag_out0[2] ),
    .X(_03224_));
 sky130_fd_sc_hd__or4_2 _05708_ (.A(_03194_),
    .B(_03196_),
    .C(_03199_),
    .D(_03224_),
    .X(_03225_));
 sky130_fd_sc_hd__or4_2 _05709_ (.A(_03219_),
    .B(_03222_),
    .C(_03223_),
    .D(_03225_),
    .X(_03226_));
 sky130_fd_sc_hd__or3_2 _05710_ (.A(_03156_),
    .B(_03158_),
    .C(_03203_),
    .X(_03227_));
 sky130_fd_sc_hd__or4b_2 _05711_ (.A(_03182_),
    .B(_03184_),
    .C(_03200_),
    .D_N(\fsm.valid0 ),
    .X(_03228_));
 sky130_fd_sc_hd__and2b_2 _05712_ (.A_N(\fsm.tag_out0[2] ),
    .B(cpu_addr[9]),
    .X(_03229_));
 sky130_fd_sc_hd__or4_2 _05713_ (.A(_03179_),
    .B(_03198_),
    .C(_03204_),
    .D(_03229_),
    .X(_03230_));
 sky130_fd_sc_hd__or3_2 _05714_ (.A(_03227_),
    .B(_03228_),
    .C(_03230_),
    .X(_03231_));
 sky130_fd_sc_hd__or4_2 _05715_ (.A(_03173_),
    .B(_03189_),
    .C(_03190_),
    .D(_03205_),
    .X(_03232_));
 sky130_fd_sc_hd__or4_2 _05716_ (.A(_03174_),
    .B(_03175_),
    .C(_03195_),
    .D(_03208_),
    .X(_03233_));
 sky130_fd_sc_hd__a2111o_2 _05717_ (.A1(_03135_),
    .A2(\fsm.tag_out0[1] ),
    .B1(_03169_),
    .C1(_03170_),
    .D1(_03185_),
    .X(_03234_));
 sky130_fd_sc_hd__or3_2 _05718_ (.A(_03232_),
    .B(_03233_),
    .C(_03234_),
    .X(_03235_));
 sky130_fd_sc_hd__nor4_2 _05719_ (.A(_03217_),
    .B(_03226_),
    .C(_03231_),
    .D(_03235_),
    .Y(_03236_));
 sky130_fd_sc_hd__xor2_2 _05720_ (.A(cpu_addr[21]),
    .B(\fsm.tag_out1[14] ),
    .X(_03237_));
 sky130_fd_sc_hd__xor2_2 _05721_ (.A(cpu_addr[29]),
    .B(\fsm.tag_out1[22] ),
    .X(_03238_));
 sky130_fd_sc_hd__xor2_2 _05722_ (.A(cpu_addr[9]),
    .B(\fsm.tag_out1[2] ),
    .X(_03239_));
 sky130_fd_sc_hd__xor2_2 _05723_ (.A(cpu_addr[11]),
    .B(\fsm.tag_out1[4] ),
    .X(_03240_));
 sky130_fd_sc_hd__or4_2 _05724_ (.A(_03237_),
    .B(_03238_),
    .C(_03239_),
    .D(_03240_),
    .X(_03241_));
 sky130_fd_sc_hd__xnor2_2 _05725_ (.A(cpu_addr[18]),
    .B(\fsm.tag_out1[11] ),
    .Y(_03242_));
 sky130_fd_sc_hd__nand2b_2 _05726_ (.A_N(cpu_addr[25]),
    .B(\fsm.tag_out1[18] ),
    .Y(_03243_));
 sky130_fd_sc_hd__and3_2 _05727_ (.A(\fsm.valid1 ),
    .B(_03242_),
    .C(_03243_),
    .X(_03244_));
 sky130_fd_sc_hd__xor2_2 _05728_ (.A(cpu_addr[26]),
    .B(\fsm.tag_out1[19] ),
    .X(_03245_));
 sky130_fd_sc_hd__xor2_2 _05729_ (.A(cpu_addr[10]),
    .B(\fsm.tag_out1[3] ),
    .X(_03246_));
 sky130_fd_sc_hd__xor2_2 _05730_ (.A(cpu_addr[15]),
    .B(\fsm.tag_out1[8] ),
    .X(_03247_));
 sky130_fd_sc_hd__and2b_2 _05731_ (.A_N(\fsm.tag_out1[9] ),
    .B(cpu_addr[16]),
    .X(_03248_));
 sky130_fd_sc_hd__and2b_2 _05732_ (.A_N(\fsm.tag_out1[12] ),
    .B(cpu_addr[19]),
    .X(_03249_));
 sky130_fd_sc_hd__and2b_2 _05733_ (.A_N(cpu_addr[14]),
    .B(\fsm.tag_out1[7] ),
    .X(_03250_));
 sky130_fd_sc_hd__and2b_2 _05734_ (.A_N(cpu_addr[28]),
    .B(\fsm.tag_out1[21] ),
    .X(_03251_));
 sky130_fd_sc_hd__and2b_2 _05735_ (.A_N(cpu_addr[22]),
    .B(\fsm.tag_out1[15] ),
    .X(_03252_));
 sky130_fd_sc_hd__or4_2 _05736_ (.A(_03249_),
    .B(_03250_),
    .C(_03251_),
    .D(_03252_),
    .X(_03253_));
 sky130_fd_sc_hd__a2111o_2 _05737_ (.A1(_03143_),
    .A2(\fsm.tag_out1[20] ),
    .B1(_03247_),
    .C1(_03248_),
    .D1(_03253_),
    .X(_03254_));
 sky130_fd_sc_hd__or4b_2 _05738_ (.A(_03245_),
    .B(_03246_),
    .C(_03254_),
    .D_N(_03244_),
    .X(_03255_));
 sky130_fd_sc_hd__a22o_2 _05739_ (.A1(cpu_addr[13]),
    .A2(_03138_),
    .B1(cpu_addr[22]),
    .B2(_03141_),
    .X(_03256_));
 sky130_fd_sc_hd__and2b_2 _05740_ (.A_N(cpu_addr[13]),
    .B(\fsm.tag_out1[6] ),
    .X(_03257_));
 sky130_fd_sc_hd__and2b_2 _05741_ (.A_N(\fsm.tag_out1[1] ),
    .B(cpu_addr[8]),
    .X(_03258_));
 sky130_fd_sc_hd__and2b_2 _05742_ (.A_N(cpu_addr[20]),
    .B(\fsm.tag_out1[13] ),
    .X(_03259_));
 sky130_fd_sc_hd__and2b_2 _05743_ (.A_N(cpu_addr[8]),
    .B(\fsm.tag_out1[1] ),
    .X(_03260_));
 sky130_fd_sc_hd__and2b_2 _05744_ (.A_N(cpu_addr[30]),
    .B(\fsm.tag_out1[23] ),
    .X(_03261_));
 sky130_fd_sc_hd__or4_2 _05745_ (.A(_03258_),
    .B(_03259_),
    .C(_03260_),
    .D(_03261_),
    .X(_03262_));
 sky130_fd_sc_hd__and2b_2 _05746_ (.A_N(\fsm.tag_out1[21] ),
    .B(cpu_addr[28]),
    .X(_03263_));
 sky130_fd_sc_hd__and2b_2 _05747_ (.A_N(\fsm.tag_out1[7] ),
    .B(cpu_addr[14]),
    .X(_03264_));
 sky130_fd_sc_hd__and2b_2 _05748_ (.A_N(cpu_addr[17]),
    .B(\fsm.tag_out1[10] ),
    .X(_03265_));
 sky130_fd_sc_hd__and2b_2 _05749_ (.A_N(cpu_addr[19]),
    .B(\fsm.tag_out1[12] ),
    .X(_03266_));
 sky130_fd_sc_hd__or4_2 _05750_ (.A(_03263_),
    .B(_03264_),
    .C(_03265_),
    .D(_03266_),
    .X(_03267_));
 sky130_fd_sc_hd__or4_2 _05751_ (.A(_03256_),
    .B(_03257_),
    .C(_03262_),
    .D(_03267_),
    .X(_03268_));
 sky130_fd_sc_hd__xor2_2 _05752_ (.A(cpu_addr[31]),
    .B(\fsm.tag_out1[24] ),
    .X(_03269_));
 sky130_fd_sc_hd__and2b_2 _05753_ (.A_N(cpu_addr[7]),
    .B(\fsm.tag_out1[0] ),
    .X(_03270_));
 sky130_fd_sc_hd__and2b_2 _05754_ (.A_N(cpu_addr[16]),
    .B(\fsm.tag_out1[9] ),
    .X(_03271_));
 sky130_fd_sc_hd__and2b_2 _05755_ (.A_N(\fsm.tag_out1[18] ),
    .B(cpu_addr[25]),
    .X(_03272_));
 sky130_fd_sc_hd__and2b_2 _05756_ (.A_N(\fsm.tag_out1[10] ),
    .B(cpu_addr[17]),
    .X(_03273_));
 sky130_fd_sc_hd__and2b_2 _05757_ (.A_N(\fsm.tag_out1[13] ),
    .B(cpu_addr[20]),
    .X(_03274_));
 sky130_fd_sc_hd__or4_2 _05758_ (.A(_03271_),
    .B(_03272_),
    .C(_03273_),
    .D(_03274_),
    .X(_03275_));
 sky130_fd_sc_hd__a2111o_2 _05759_ (.A1(cpu_addr[27]),
    .A2(_03144_),
    .B1(_03269_),
    .C1(_03270_),
    .D1(_03275_),
    .X(_03276_));
 sky130_fd_sc_hd__and2b_2 _05760_ (.A_N(\fsm.tag_out1[17] ),
    .B(cpu_addr[24]),
    .X(_03277_));
 sky130_fd_sc_hd__and2b_2 _05761_ (.A_N(cpu_addr[24]),
    .B(\fsm.tag_out1[17] ),
    .X(_03278_));
 sky130_fd_sc_hd__and2b_2 _05762_ (.A_N(\fsm.tag_out1[0] ),
    .B(cpu_addr[7]),
    .X(_03279_));
 sky130_fd_sc_hd__and2b_2 _05763_ (.A_N(\fsm.tag_out1[23] ),
    .B(cpu_addr[30]),
    .X(_03280_));
 sky130_fd_sc_hd__or4_2 _05764_ (.A(_03277_),
    .B(_03278_),
    .C(_03279_),
    .D(_03280_),
    .X(_03281_));
 sky130_fd_sc_hd__xor2_2 _05765_ (.A(cpu_addr[12]),
    .B(\fsm.tag_out1[5] ),
    .X(_03282_));
 sky130_fd_sc_hd__xor2_2 _05766_ (.A(cpu_addr[23]),
    .B(\fsm.tag_out1[16] ),
    .X(_03283_));
 sky130_fd_sc_hd__or4_2 _05767_ (.A(_03276_),
    .B(_03281_),
    .C(_03282_),
    .D(_03283_),
    .X(_03284_));
 sky130_fd_sc_hd__or4_2 _05768_ (.A(_03241_),
    .B(_03255_),
    .C(_03268_),
    .D(_03284_),
    .X(_03285_));
 sky130_fd_sc_hd__nand2_2 _05769_ (.A(cpu_addr[27]),
    .B(\fsm.tag_out1[20] ),
    .Y(_03286_));
 sky130_fd_sc_hd__or2_2 _05770_ (.A(cpu_addr[27]),
    .B(\fsm.tag_out1[20] ),
    .X(_03287_));
 sky130_fd_sc_hd__a211o_2 _05771_ (.A1(_03286_),
    .A2(_03287_),
    .B1(_03238_),
    .C1(_03269_),
    .X(_03288_));
 sky130_fd_sc_hd__and2b_2 _05772_ (.A_N(cpu_addr[11]),
    .B(\fsm.tag_out1[4] ),
    .X(_03289_));
 sky130_fd_sc_hd__or3_2 _05773_ (.A(_03247_),
    .B(_03248_),
    .C(_03289_),
    .X(_03290_));
 sky130_fd_sc_hd__nand2_2 _05774_ (.A(cpu_addr[17]),
    .B(\fsm.tag_out1[10] ),
    .Y(_03291_));
 sky130_fd_sc_hd__or2_2 _05775_ (.A(cpu_addr[17]),
    .B(\fsm.tag_out1[10] ),
    .X(_03292_));
 sky130_fd_sc_hd__a211o_2 _05776_ (.A1(_03291_),
    .A2(_03292_),
    .B1(_03263_),
    .C1(_03266_),
    .X(_03293_));
 sky130_fd_sc_hd__or3_2 _05777_ (.A(_03288_),
    .B(_03290_),
    .C(_03293_),
    .X(_03294_));
 sky130_fd_sc_hd__or3_2 _05778_ (.A(_03259_),
    .B(_03264_),
    .C(_03274_),
    .X(_03295_));
 sky130_fd_sc_hd__and2b_2 _05779_ (.A_N(\fsm.tag_out1[4] ),
    .B(cpu_addr[11]),
    .X(_03296_));
 sky130_fd_sc_hd__or4_2 _05780_ (.A(_03249_),
    .B(_03250_),
    .C(_03260_),
    .D(_03296_),
    .X(_03297_));
 sky130_fd_sc_hd__and2b_2 _05781_ (.A_N(\fsm.tag_out1[11] ),
    .B(cpu_addr[18]),
    .X(_03298_));
 sky130_fd_sc_hd__a2111o_2 _05782_ (.A1(cpu_addr[13]),
    .A2(_03138_),
    .B1(_03271_),
    .C1(_03272_),
    .D1(_03298_),
    .X(_03299_));
 sky130_fd_sc_hd__and2b_2 _05783_ (.A_N(cpu_addr[18]),
    .B(\fsm.tag_out1[11] ),
    .X(_03300_));
 sky130_fd_sc_hd__and2b_2 _05784_ (.A_N(cpu_addr[10]),
    .B(\fsm.tag_out1[3] ),
    .X(_03301_));
 sky130_fd_sc_hd__a2111o_2 _05785_ (.A1(cpu_addr[22]),
    .A2(_03141_),
    .B1(_03257_),
    .C1(_03300_),
    .D1(_03301_),
    .X(_03302_));
 sky130_fd_sc_hd__or4_2 _05786_ (.A(_03295_),
    .B(_03297_),
    .C(_03299_),
    .D(_03302_),
    .X(_03303_));
 sky130_fd_sc_hd__o21ai_2 _05787_ (.A1(_03136_),
    .A2(\fsm.tag_out1[2] ),
    .B1(\fsm.valid1 ),
    .Y(_03304_));
 sky130_fd_sc_hd__a21o_2 _05788_ (.A1(_03136_),
    .A2(\fsm.tag_out1[2] ),
    .B1(_03277_),
    .X(_03305_));
 sky130_fd_sc_hd__or4_2 _05789_ (.A(_03251_),
    .B(_03258_),
    .C(_03270_),
    .D(_03278_),
    .X(_03306_));
 sky130_fd_sc_hd__or4_2 _05790_ (.A(_03283_),
    .B(_03304_),
    .C(_03305_),
    .D(_03306_),
    .X(_03307_));
 sky130_fd_sc_hd__and2b_2 _05791_ (.A_N(cpu_addr[26]),
    .B(\fsm.tag_out1[19] ),
    .X(_03308_));
 sky130_fd_sc_hd__a2111o_2 _05792_ (.A1(cpu_addr[10]),
    .A2(_03137_),
    .B1(_03252_),
    .C1(_03261_),
    .D1(_03308_),
    .X(_03309_));
 sky130_fd_sc_hd__a21o_2 _05793_ (.A1(_03140_),
    .A2(\fsm.tag_out1[14] ),
    .B1(_03279_),
    .X(_03310_));
 sky130_fd_sc_hd__o21ai_2 _05794_ (.A1(_03140_),
    .A2(\fsm.tag_out1[14] ),
    .B1(_03243_),
    .Y(_03311_));
 sky130_fd_sc_hd__and2b_2 _05795_ (.A_N(\fsm.tag_out1[19] ),
    .B(cpu_addr[26]),
    .X(_03312_));
 sky130_fd_sc_hd__or3_2 _05796_ (.A(_03280_),
    .B(_03282_),
    .C(_03312_),
    .X(_03313_));
 sky130_fd_sc_hd__or4_2 _05797_ (.A(_03309_),
    .B(_03310_),
    .C(_03311_),
    .D(_03313_),
    .X(_03314_));
 sky130_fd_sc_hd__nor4_2 _05798_ (.A(_03294_),
    .B(_03303_),
    .C(_03307_),
    .D(_03314_),
    .Y(_03315_));
 sky130_fd_sc_hd__or4_2 _05799_ (.A(_03182_),
    .B(_03184_),
    .C(_03200_),
    .D(_03209_),
    .X(_03316_));
 sky130_fd_sc_hd__or2_2 _05800_ (.A(_03155_),
    .B(_03157_),
    .X(_03317_));
 sky130_fd_sc_hd__or4_2 _05801_ (.A(_03178_),
    .B(_03179_),
    .C(_03198_),
    .D(_03229_),
    .X(_03318_));
 sky130_fd_sc_hd__or4_2 _05802_ (.A(_03172_),
    .B(_03183_),
    .C(_03204_),
    .D(_03207_),
    .X(_03319_));
 sky130_fd_sc_hd__or4_2 _05803_ (.A(_03316_),
    .B(_03317_),
    .C(_03318_),
    .D(_03319_),
    .X(_03320_));
 sky130_fd_sc_hd__or2_2 _05804_ (.A(_03195_),
    .B(_03201_),
    .X(_03321_));
 sky130_fd_sc_hd__and2b_2 _05805_ (.A_N(\fsm.tag_out0[23] ),
    .B(cpu_addr[30]),
    .X(_03322_));
 sky130_fd_sc_hd__and2b_2 _05806_ (.A_N(cpu_addr[30]),
    .B(\fsm.tag_out0[23] ),
    .X(_03323_));
 sky130_fd_sc_hd__or4_2 _05807_ (.A(_03174_),
    .B(_03175_),
    .C(_03322_),
    .D(_03323_),
    .X(_03324_));
 sky130_fd_sc_hd__or4_2 _05808_ (.A(_03169_),
    .B(_03185_),
    .C(_03208_),
    .D(_03224_),
    .X(_03325_));
 sky130_fd_sc_hd__or4_2 _05809_ (.A(_03199_),
    .B(_03321_),
    .C(_03324_),
    .D(_03325_),
    .X(_03326_));
 sky130_fd_sc_hd__or4_2 _05810_ (.A(_03156_),
    .B(_03158_),
    .C(_03203_),
    .D(_03214_),
    .X(_03327_));
 sky130_fd_sc_hd__a2111o_2 _05811_ (.A1(_03135_),
    .A2(\fsm.tag_out0[1] ),
    .B1(_03170_),
    .C1(_03194_),
    .D1(_03196_),
    .X(_03328_));
 sky130_fd_sc_hd__or4_2 _05812_ (.A(_03180_),
    .B(_03189_),
    .C(_03205_),
    .D(_03210_),
    .X(_03329_));
 sky130_fd_sc_hd__or4b_2 _05813_ (.A(_03160_),
    .B(_03168_),
    .C(_03190_),
    .D_N(\fsm.valid0 ),
    .X(_03330_));
 sky130_fd_sc_hd__or4_2 _05814_ (.A(_03173_),
    .B(_03187_),
    .C(_03188_),
    .D(_03218_),
    .X(_03331_));
 sky130_fd_sc_hd__or4_2 _05815_ (.A(_03328_),
    .B(_03329_),
    .C(_03330_),
    .D(_03331_),
    .X(_03332_));
 sky130_fd_sc_hd__nor4_2 _05816_ (.A(_03320_),
    .B(_03326_),
    .C(_03327_),
    .D(_03332_),
    .Y(_03333_));
 sky130_fd_sc_hd__or3_2 _05817_ (.A(_03239_),
    .B(_03277_),
    .C(_03289_),
    .X(_03334_));
 sky130_fd_sc_hd__or4_2 _05818_ (.A(_03248_),
    .B(_03265_),
    .C(_03273_),
    .D(_03278_),
    .X(_03335_));
 sky130_fd_sc_hd__or4_2 _05819_ (.A(_03251_),
    .B(_03263_),
    .C(_03266_),
    .D(_03270_),
    .X(_03336_));
 sky130_fd_sc_hd__or4_2 _05820_ (.A(_03258_),
    .B(_03271_),
    .C(_03272_),
    .D(_03279_),
    .X(_03337_));
 sky130_fd_sc_hd__or4_2 _05821_ (.A(_03334_),
    .B(_03335_),
    .C(_03336_),
    .D(_03337_),
    .X(_03338_));
 sky130_fd_sc_hd__o21ai_2 _05822_ (.A1(_03139_),
    .A2(\fsm.tag_out1[11] ),
    .B1(_03243_),
    .Y(_03339_));
 sky130_fd_sc_hd__or4_2 _05823_ (.A(_03280_),
    .B(_03282_),
    .C(_03301_),
    .D(_03312_),
    .X(_03340_));
 sky130_fd_sc_hd__or4_2 _05824_ (.A(_03237_),
    .B(_03256_),
    .C(_03339_),
    .D(_03340_),
    .X(_03341_));
 sky130_fd_sc_hd__or2_2 _05825_ (.A(_03247_),
    .B(_03288_),
    .X(_03342_));
 sky130_fd_sc_hd__or4_2 _05826_ (.A(_03257_),
    .B(_03260_),
    .C(_03296_),
    .D(_03300_),
    .X(_03343_));
 sky130_fd_sc_hd__or4_2 _05827_ (.A(_03249_),
    .B(_03250_),
    .C(_03259_),
    .D(_03264_),
    .X(_03344_));
 sky130_fd_sc_hd__or3b_2 _05828_ (.A(_03274_),
    .B(_03283_),
    .C_N(\fsm.valid1 ),
    .X(_03345_));
 sky130_fd_sc_hd__or4_2 _05829_ (.A(_03309_),
    .B(_03343_),
    .C(_03344_),
    .D(_03345_),
    .X(_03346_));
 sky130_fd_sc_hd__nor4_2 _05830_ (.A(_03338_),
    .B(_03341_),
    .C(_03342_),
    .D(_03346_),
    .Y(_03347_));
 sky130_fd_sc_hd__and2_2 _05831_ (.A(\data_array.rdata1[0] ),
    .B(_03347_),
    .X(_03348_));
 sky130_fd_sc_hd__mux2_1 _05832_ (.A0(_03348_),
    .A1(\data_array.rdata0[0] ),
    .S(_03333_),
    .X(_03349_));
 sky130_fd_sc_hd__a22o_2 _05833_ (.A1(mem_rdata[0]),
    .A2(_03153_),
    .B1(_03154_),
    .B2(_03349_),
    .X(cpu_rdata[0]));
 sky130_fd_sc_hd__o21a_2 _05834_ (.A1(\data_array.rdata0[1] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03350_));
 sky130_fd_sc_hd__a21o_2 _05835_ (.A1(\data_array.rdata1[1] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03351_));
 sky130_fd_sc_hd__a22o_2 _05836_ (.A1(mem_rdata[1]),
    .A2(_03153_),
    .B1(_03350_),
    .B2(_03351_),
    .X(cpu_rdata[1]));
 sky130_fd_sc_hd__o21a_2 _05837_ (.A1(\data_array.rdata0[2] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03352_));
 sky130_fd_sc_hd__a21o_2 _05838_ (.A1(\data_array.rdata1[2] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03353_));
 sky130_fd_sc_hd__a22o_2 _05839_ (.A1(mem_rdata[2]),
    .A2(_03153_),
    .B1(_03352_),
    .B2(_03353_),
    .X(cpu_rdata[2]));
 sky130_fd_sc_hd__o21a_2 _05840_ (.A1(\data_array.rdata0[3] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03354_));
 sky130_fd_sc_hd__a21o_2 _05841_ (.A1(\data_array.rdata1[3] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03355_));
 sky130_fd_sc_hd__a22o_2 _05842_ (.A1(mem_rdata[3]),
    .A2(_03153_),
    .B1(_03354_),
    .B2(_03355_),
    .X(cpu_rdata[3]));
 sky130_fd_sc_hd__o21a_2 _05843_ (.A1(\data_array.rdata0[4] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03356_));
 sky130_fd_sc_hd__a21o_2 _05844_ (.A1(\data_array.rdata1[4] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03357_));
 sky130_fd_sc_hd__a22o_2 _05845_ (.A1(mem_rdata[4]),
    .A2(_03153_),
    .B1(_03356_),
    .B2(_03357_),
    .X(cpu_rdata[4]));
 sky130_fd_sc_hd__o21a_2 _05846_ (.A1(\data_array.rdata0[5] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03358_));
 sky130_fd_sc_hd__a21o_2 _05847_ (.A1(\data_array.rdata1[5] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03359_));
 sky130_fd_sc_hd__a22o_2 _05848_ (.A1(mem_rdata[5]),
    .A2(_03153_),
    .B1(_03358_),
    .B2(_03359_),
    .X(cpu_rdata[5]));
 sky130_fd_sc_hd__o21a_2 _05849_ (.A1(\data_array.rdata0[6] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03360_));
 sky130_fd_sc_hd__a21o_2 _05850_ (.A1(\data_array.rdata1[6] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03361_));
 sky130_fd_sc_hd__a22o_2 _05851_ (.A1(mem_rdata[6]),
    .A2(_03153_),
    .B1(_03360_),
    .B2(_03361_),
    .X(cpu_rdata[6]));
 sky130_fd_sc_hd__o21a_2 _05852_ (.A1(\data_array.rdata0[7] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03362_));
 sky130_fd_sc_hd__a21o_2 _05853_ (.A1(\data_array.rdata1[7] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03363_));
 sky130_fd_sc_hd__a22o_2 _05854_ (.A1(mem_rdata[7]),
    .A2(_03153_),
    .B1(_03362_),
    .B2(_03363_),
    .X(cpu_rdata[7]));
 sky130_fd_sc_hd__o21a_2 _05855_ (.A1(\data_array.rdata0[8] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03364_));
 sky130_fd_sc_hd__a21o_2 _05856_ (.A1(\data_array.rdata1[8] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03365_));
 sky130_fd_sc_hd__a22o_2 _05857_ (.A1(mem_rdata[8]),
    .A2(_03153_),
    .B1(_03364_),
    .B2(_03365_),
    .X(cpu_rdata[8]));
 sky130_fd_sc_hd__o21a_2 _05858_ (.A1(\data_array.rdata0[9] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03366_));
 sky130_fd_sc_hd__a21o_2 _05859_ (.A1(\data_array.rdata1[9] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03367_));
 sky130_fd_sc_hd__a22o_2 _05860_ (.A1(mem_rdata[9]),
    .A2(_03153_),
    .B1(_03366_),
    .B2(_03367_),
    .X(cpu_rdata[9]));
 sky130_fd_sc_hd__o21a_2 _05861_ (.A1(\data_array.rdata0[10] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03368_));
 sky130_fd_sc_hd__a21o_2 _05862_ (.A1(\data_array.rdata1[10] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03369_));
 sky130_fd_sc_hd__a22o_2 _05863_ (.A1(mem_rdata[10]),
    .A2(_03153_),
    .B1(_03368_),
    .B2(_03369_),
    .X(cpu_rdata[10]));
 sky130_fd_sc_hd__o21a_2 _05864_ (.A1(\data_array.rdata0[11] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03370_));
 sky130_fd_sc_hd__a21o_2 _05865_ (.A1(\data_array.rdata1[11] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03371_));
 sky130_fd_sc_hd__a22o_2 _05866_ (.A1(mem_rdata[11]),
    .A2(_03153_),
    .B1(_03370_),
    .B2(_03371_),
    .X(cpu_rdata[11]));
 sky130_fd_sc_hd__o21a_2 _05867_ (.A1(\data_array.rdata0[12] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03372_));
 sky130_fd_sc_hd__a21o_2 _05868_ (.A1(\data_array.rdata1[12] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03373_));
 sky130_fd_sc_hd__a22o_2 _05869_ (.A1(mem_rdata[12]),
    .A2(_03153_),
    .B1(_03372_),
    .B2(_03373_),
    .X(cpu_rdata[12]));
 sky130_fd_sc_hd__o21a_2 _05870_ (.A1(\data_array.rdata0[13] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03374_));
 sky130_fd_sc_hd__a21o_2 _05871_ (.A1(\data_array.rdata1[13] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03375_));
 sky130_fd_sc_hd__a22o_2 _05872_ (.A1(mem_rdata[13]),
    .A2(_03153_),
    .B1(_03374_),
    .B2(_03375_),
    .X(cpu_rdata[13]));
 sky130_fd_sc_hd__o21a_2 _05873_ (.A1(\data_array.rdata0[14] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03376_));
 sky130_fd_sc_hd__a21o_2 _05874_ (.A1(\data_array.rdata1[14] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03377_));
 sky130_fd_sc_hd__a22o_2 _05875_ (.A1(mem_rdata[14]),
    .A2(_03153_),
    .B1(_03376_),
    .B2(_03377_),
    .X(cpu_rdata[14]));
 sky130_fd_sc_hd__o21a_2 _05876_ (.A1(\data_array.rdata0[15] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03378_));
 sky130_fd_sc_hd__a21o_2 _05877_ (.A1(\data_array.rdata1[15] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03379_));
 sky130_fd_sc_hd__a22o_2 _05878_ (.A1(mem_rdata[15]),
    .A2(_03153_),
    .B1(_03378_),
    .B2(_03379_),
    .X(cpu_rdata[15]));
 sky130_fd_sc_hd__o21a_2 _05879_ (.A1(\data_array.rdata0[16] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03380_));
 sky130_fd_sc_hd__a21o_2 _05880_ (.A1(\data_array.rdata1[16] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03381_));
 sky130_fd_sc_hd__a22o_2 _05881_ (.A1(mem_rdata[16]),
    .A2(_03153_),
    .B1(_03380_),
    .B2(_03381_),
    .X(cpu_rdata[16]));
 sky130_fd_sc_hd__o21a_2 _05882_ (.A1(\data_array.rdata0[17] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03382_));
 sky130_fd_sc_hd__a21o_2 _05883_ (.A1(\data_array.rdata1[17] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03383_));
 sky130_fd_sc_hd__a22o_2 _05884_ (.A1(mem_rdata[17]),
    .A2(_03153_),
    .B1(_03382_),
    .B2(_03383_),
    .X(cpu_rdata[17]));
 sky130_fd_sc_hd__o21a_2 _05885_ (.A1(\data_array.rdata0[18] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03384_));
 sky130_fd_sc_hd__a21o_2 _05886_ (.A1(\data_array.rdata1[18] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03385_));
 sky130_fd_sc_hd__a22o_2 _05887_ (.A1(mem_rdata[18]),
    .A2(_03153_),
    .B1(_03384_),
    .B2(_03385_),
    .X(cpu_rdata[18]));
 sky130_fd_sc_hd__o21a_2 _05888_ (.A1(\data_array.rdata0[19] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03386_));
 sky130_fd_sc_hd__a21o_2 _05889_ (.A1(\data_array.rdata1[19] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03387_));
 sky130_fd_sc_hd__a22o_2 _05890_ (.A1(mem_rdata[19]),
    .A2(_03153_),
    .B1(_03386_),
    .B2(_03387_),
    .X(cpu_rdata[19]));
 sky130_fd_sc_hd__o21a_2 _05891_ (.A1(\data_array.rdata0[20] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03388_));
 sky130_fd_sc_hd__a21o_2 _05892_ (.A1(\data_array.rdata1[20] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03389_));
 sky130_fd_sc_hd__a22o_2 _05893_ (.A1(mem_rdata[20]),
    .A2(_03153_),
    .B1(_03388_),
    .B2(_03389_),
    .X(cpu_rdata[20]));
 sky130_fd_sc_hd__o21a_2 _05894_ (.A1(\data_array.rdata0[21] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03390_));
 sky130_fd_sc_hd__a21o_2 _05895_ (.A1(\data_array.rdata1[21] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03391_));
 sky130_fd_sc_hd__a22o_2 _05896_ (.A1(mem_rdata[21]),
    .A2(_03153_),
    .B1(_03390_),
    .B2(_03391_),
    .X(cpu_rdata[21]));
 sky130_fd_sc_hd__o21a_2 _05897_ (.A1(\data_array.rdata0[22] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03392_));
 sky130_fd_sc_hd__a21o_2 _05898_ (.A1(\data_array.rdata1[22] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03393_));
 sky130_fd_sc_hd__a22o_2 _05899_ (.A1(mem_rdata[22]),
    .A2(_03153_),
    .B1(_03392_),
    .B2(_03393_),
    .X(cpu_rdata[22]));
 sky130_fd_sc_hd__o21a_2 _05900_ (.A1(\data_array.rdata0[23] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03394_));
 sky130_fd_sc_hd__a21o_2 _05901_ (.A1(\data_array.rdata1[23] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03395_));
 sky130_fd_sc_hd__a22o_2 _05902_ (.A1(mem_rdata[23]),
    .A2(_03153_),
    .B1(_03394_),
    .B2(_03395_),
    .X(cpu_rdata[23]));
 sky130_fd_sc_hd__o21a_2 _05903_ (.A1(\data_array.rdata0[24] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03396_));
 sky130_fd_sc_hd__a21o_2 _05904_ (.A1(\data_array.rdata1[24] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03397_));
 sky130_fd_sc_hd__a22o_2 _05905_ (.A1(mem_rdata[24]),
    .A2(_03153_),
    .B1(_03396_),
    .B2(_03397_),
    .X(cpu_rdata[24]));
 sky130_fd_sc_hd__o21a_2 _05906_ (.A1(\data_array.rdata0[25] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03398_));
 sky130_fd_sc_hd__a21o_2 _05907_ (.A1(\data_array.rdata1[25] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03399_));
 sky130_fd_sc_hd__a22o_2 _05908_ (.A1(mem_rdata[25]),
    .A2(_03153_),
    .B1(_03398_),
    .B2(_03399_),
    .X(cpu_rdata[25]));
 sky130_fd_sc_hd__o21a_2 _05909_ (.A1(\data_array.rdata0[26] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03400_));
 sky130_fd_sc_hd__a21o_2 _05910_ (.A1(\data_array.rdata1[26] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03401_));
 sky130_fd_sc_hd__a22o_2 _05911_ (.A1(mem_rdata[26]),
    .A2(_03153_),
    .B1(_03400_),
    .B2(_03401_),
    .X(cpu_rdata[26]));
 sky130_fd_sc_hd__o21a_2 _05912_ (.A1(\data_array.rdata0[27] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03402_));
 sky130_fd_sc_hd__a21o_2 _05913_ (.A1(\data_array.rdata1[27] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03403_));
 sky130_fd_sc_hd__a22o_2 _05914_ (.A1(mem_rdata[27]),
    .A2(_03153_),
    .B1(_03402_),
    .B2(_03403_),
    .X(cpu_rdata[27]));
 sky130_fd_sc_hd__o21a_2 _05915_ (.A1(\data_array.rdata0[28] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03404_));
 sky130_fd_sc_hd__a21o_2 _05916_ (.A1(\data_array.rdata1[28] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03405_));
 sky130_fd_sc_hd__a22o_2 _05917_ (.A1(mem_rdata[28]),
    .A2(_03153_),
    .B1(_03404_),
    .B2(_03405_),
    .X(cpu_rdata[28]));
 sky130_fd_sc_hd__o21a_2 _05918_ (.A1(\data_array.rdata0[29] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03406_));
 sky130_fd_sc_hd__a21o_2 _05919_ (.A1(\data_array.rdata1[29] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03407_));
 sky130_fd_sc_hd__a22o_2 _05920_ (.A1(mem_rdata[29]),
    .A2(_03153_),
    .B1(_03406_),
    .B2(_03407_),
    .X(cpu_rdata[29]));
 sky130_fd_sc_hd__o21a_2 _05921_ (.A1(\data_array.rdata0[30] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03408_));
 sky130_fd_sc_hd__a21o_2 _05922_ (.A1(\data_array.rdata1[30] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03409_));
 sky130_fd_sc_hd__a22o_2 _05923_ (.A1(mem_rdata[30]),
    .A2(_03153_),
    .B1(_03408_),
    .B2(_03409_),
    .X(cpu_rdata[30]));
 sky130_fd_sc_hd__o21a_2 _05924_ (.A1(\data_array.rdata0[31] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03410_));
 sky130_fd_sc_hd__a21o_2 _05925_ (.A1(\data_array.rdata1[31] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03411_));
 sky130_fd_sc_hd__a22o_2 _05926_ (.A1(mem_rdata[31]),
    .A2(_03153_),
    .B1(_03410_),
    .B2(_03411_),
    .X(cpu_rdata[31]));
 sky130_fd_sc_hd__o21a_2 _05927_ (.A1(\data_array.rdata0[32] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03412_));
 sky130_fd_sc_hd__a21o_2 _05928_ (.A1(\data_array.rdata1[32] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03413_));
 sky130_fd_sc_hd__a22o_2 _05929_ (.A1(mem_rdata[32]),
    .A2(_03153_),
    .B1(_03412_),
    .B2(_03413_),
    .X(cpu_rdata[32]));
 sky130_fd_sc_hd__o21a_2 _05930_ (.A1(\data_array.rdata0[33] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03414_));
 sky130_fd_sc_hd__a21o_2 _05931_ (.A1(\data_array.rdata1[33] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03415_));
 sky130_fd_sc_hd__a22o_2 _05932_ (.A1(mem_rdata[33]),
    .A2(_03153_),
    .B1(_03414_),
    .B2(_03415_),
    .X(cpu_rdata[33]));
 sky130_fd_sc_hd__o21a_2 _05933_ (.A1(\data_array.rdata0[34] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03416_));
 sky130_fd_sc_hd__a21o_2 _05934_ (.A1(\data_array.rdata1[34] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03417_));
 sky130_fd_sc_hd__a22o_2 _05935_ (.A1(mem_rdata[34]),
    .A2(_03153_),
    .B1(_03416_),
    .B2(_03417_),
    .X(cpu_rdata[34]));
 sky130_fd_sc_hd__o21a_2 _05936_ (.A1(\data_array.rdata0[35] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03418_));
 sky130_fd_sc_hd__a21o_2 _05937_ (.A1(\data_array.rdata1[35] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03419_));
 sky130_fd_sc_hd__a22o_2 _05938_ (.A1(mem_rdata[35]),
    .A2(_03153_),
    .B1(_03418_),
    .B2(_03419_),
    .X(cpu_rdata[35]));
 sky130_fd_sc_hd__o21a_2 _05939_ (.A1(\data_array.rdata0[36] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03420_));
 sky130_fd_sc_hd__a21o_2 _05940_ (.A1(\data_array.rdata1[36] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03421_));
 sky130_fd_sc_hd__a22o_2 _05941_ (.A1(mem_rdata[36]),
    .A2(_03153_),
    .B1(_03420_),
    .B2(_03421_),
    .X(cpu_rdata[36]));
 sky130_fd_sc_hd__o21a_2 _05942_ (.A1(\data_array.rdata0[37] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03422_));
 sky130_fd_sc_hd__a21o_2 _05943_ (.A1(\data_array.rdata1[37] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03423_));
 sky130_fd_sc_hd__a22o_2 _05944_ (.A1(mem_rdata[37]),
    .A2(_03153_),
    .B1(_03422_),
    .B2(_03423_),
    .X(cpu_rdata[37]));
 sky130_fd_sc_hd__o21a_2 _05945_ (.A1(\data_array.rdata0[38] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03424_));
 sky130_fd_sc_hd__a21o_2 _05946_ (.A1(\data_array.rdata1[38] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03425_));
 sky130_fd_sc_hd__a22o_2 _05947_ (.A1(mem_rdata[38]),
    .A2(_03153_),
    .B1(_03424_),
    .B2(_03425_),
    .X(cpu_rdata[38]));
 sky130_fd_sc_hd__o21a_2 _05948_ (.A1(\data_array.rdata0[39] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03426_));
 sky130_fd_sc_hd__a21o_2 _05949_ (.A1(\data_array.rdata1[39] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03427_));
 sky130_fd_sc_hd__a22o_2 _05950_ (.A1(mem_rdata[39]),
    .A2(_03153_),
    .B1(_03426_),
    .B2(_03427_),
    .X(cpu_rdata[39]));
 sky130_fd_sc_hd__o21a_2 _05951_ (.A1(\data_array.rdata0[40] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03428_));
 sky130_fd_sc_hd__a21o_2 _05952_ (.A1(\data_array.rdata1[40] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03429_));
 sky130_fd_sc_hd__a22o_2 _05953_ (.A1(mem_rdata[40]),
    .A2(_03153_),
    .B1(_03428_),
    .B2(_03429_),
    .X(cpu_rdata[40]));
 sky130_fd_sc_hd__o21a_2 _05954_ (.A1(\data_array.rdata0[41] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03430_));
 sky130_fd_sc_hd__a21o_2 _05955_ (.A1(\data_array.rdata1[41] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03431_));
 sky130_fd_sc_hd__a22o_2 _05956_ (.A1(mem_rdata[41]),
    .A2(_03153_),
    .B1(_03430_),
    .B2(_03431_),
    .X(cpu_rdata[41]));
 sky130_fd_sc_hd__o21a_2 _05957_ (.A1(\data_array.rdata0[42] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03432_));
 sky130_fd_sc_hd__a21o_2 _05958_ (.A1(\data_array.rdata1[42] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03433_));
 sky130_fd_sc_hd__a22o_2 _05959_ (.A1(mem_rdata[42]),
    .A2(_03153_),
    .B1(_03432_),
    .B2(_03433_),
    .X(cpu_rdata[42]));
 sky130_fd_sc_hd__o21a_2 _05960_ (.A1(\data_array.rdata0[43] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03434_));
 sky130_fd_sc_hd__a21o_2 _05961_ (.A1(\data_array.rdata1[43] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03435_));
 sky130_fd_sc_hd__a22o_2 _05962_ (.A1(mem_rdata[43]),
    .A2(_03153_),
    .B1(_03434_),
    .B2(_03435_),
    .X(cpu_rdata[43]));
 sky130_fd_sc_hd__o21a_2 _05963_ (.A1(\data_array.rdata0[44] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03436_));
 sky130_fd_sc_hd__a21o_2 _05964_ (.A1(\data_array.rdata1[44] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03437_));
 sky130_fd_sc_hd__a22o_2 _05965_ (.A1(mem_rdata[44]),
    .A2(_03153_),
    .B1(_03436_),
    .B2(_03437_),
    .X(cpu_rdata[44]));
 sky130_fd_sc_hd__o21a_2 _05966_ (.A1(\data_array.rdata0[45] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03438_));
 sky130_fd_sc_hd__a21o_2 _05967_ (.A1(\data_array.rdata1[45] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03439_));
 sky130_fd_sc_hd__a22o_2 _05968_ (.A1(mem_rdata[45]),
    .A2(_03153_),
    .B1(_03438_),
    .B2(_03439_),
    .X(cpu_rdata[45]));
 sky130_fd_sc_hd__o21a_2 _05969_ (.A1(\data_array.rdata0[46] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03440_));
 sky130_fd_sc_hd__a21o_2 _05970_ (.A1(\data_array.rdata1[46] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03441_));
 sky130_fd_sc_hd__a22o_2 _05971_ (.A1(mem_rdata[46]),
    .A2(_03153_),
    .B1(_03440_),
    .B2(_03441_),
    .X(cpu_rdata[46]));
 sky130_fd_sc_hd__o21a_2 _05972_ (.A1(\data_array.rdata0[47] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03442_));
 sky130_fd_sc_hd__a21o_2 _05973_ (.A1(\data_array.rdata1[47] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03443_));
 sky130_fd_sc_hd__a22o_2 _05974_ (.A1(mem_rdata[47]),
    .A2(_03153_),
    .B1(_03442_),
    .B2(_03443_),
    .X(cpu_rdata[47]));
 sky130_fd_sc_hd__o21a_2 _05975_ (.A1(\data_array.rdata0[48] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03444_));
 sky130_fd_sc_hd__a21o_2 _05976_ (.A1(\data_array.rdata1[48] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03445_));
 sky130_fd_sc_hd__a22o_2 _05977_ (.A1(mem_rdata[48]),
    .A2(_03153_),
    .B1(_03444_),
    .B2(_03445_),
    .X(cpu_rdata[48]));
 sky130_fd_sc_hd__o21a_2 _05978_ (.A1(\data_array.rdata0[49] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03446_));
 sky130_fd_sc_hd__a21o_2 _05979_ (.A1(\data_array.rdata1[49] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03447_));
 sky130_fd_sc_hd__a22o_2 _05980_ (.A1(mem_rdata[49]),
    .A2(_03153_),
    .B1(_03446_),
    .B2(_03447_),
    .X(cpu_rdata[49]));
 sky130_fd_sc_hd__o21a_2 _05981_ (.A1(\data_array.rdata0[50] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03448_));
 sky130_fd_sc_hd__a21o_2 _05982_ (.A1(\data_array.rdata1[50] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03449_));
 sky130_fd_sc_hd__a22o_2 _05983_ (.A1(mem_rdata[50]),
    .A2(_03153_),
    .B1(_03448_),
    .B2(_03449_),
    .X(cpu_rdata[50]));
 sky130_fd_sc_hd__o21a_2 _05984_ (.A1(\data_array.rdata0[51] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03450_));
 sky130_fd_sc_hd__a21o_2 _05985_ (.A1(\data_array.rdata1[51] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03451_));
 sky130_fd_sc_hd__a22o_2 _05986_ (.A1(mem_rdata[51]),
    .A2(_03153_),
    .B1(_03450_),
    .B2(_03451_),
    .X(cpu_rdata[51]));
 sky130_fd_sc_hd__o21a_2 _05987_ (.A1(\data_array.rdata0[52] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03452_));
 sky130_fd_sc_hd__a21o_2 _05988_ (.A1(\data_array.rdata1[52] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03453_));
 sky130_fd_sc_hd__a22o_2 _05989_ (.A1(mem_rdata[52]),
    .A2(_03153_),
    .B1(_03452_),
    .B2(_03453_),
    .X(cpu_rdata[52]));
 sky130_fd_sc_hd__o21a_2 _05990_ (.A1(\data_array.rdata0[53] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03454_));
 sky130_fd_sc_hd__a21o_2 _05991_ (.A1(\data_array.rdata1[53] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03455_));
 sky130_fd_sc_hd__a22o_2 _05992_ (.A1(mem_rdata[53]),
    .A2(_03153_),
    .B1(_03454_),
    .B2(_03455_),
    .X(cpu_rdata[53]));
 sky130_fd_sc_hd__o21a_2 _05993_ (.A1(\data_array.rdata0[54] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03456_));
 sky130_fd_sc_hd__a21o_2 _05994_ (.A1(\data_array.rdata1[54] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03457_));
 sky130_fd_sc_hd__a22o_2 _05995_ (.A1(mem_rdata[54]),
    .A2(_03153_),
    .B1(_03456_),
    .B2(_03457_),
    .X(cpu_rdata[54]));
 sky130_fd_sc_hd__o21a_2 _05996_ (.A1(\data_array.rdata0[55] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03458_));
 sky130_fd_sc_hd__a21o_2 _05997_ (.A1(\data_array.rdata1[55] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03459_));
 sky130_fd_sc_hd__a22o_2 _05998_ (.A1(mem_rdata[55]),
    .A2(_03153_),
    .B1(_03458_),
    .B2(_03459_),
    .X(cpu_rdata[55]));
 sky130_fd_sc_hd__o21a_2 _05999_ (.A1(\data_array.rdata0[56] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03460_));
 sky130_fd_sc_hd__a21o_2 _06000_ (.A1(\data_array.rdata1[56] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03461_));
 sky130_fd_sc_hd__a22o_2 _06001_ (.A1(mem_rdata[56]),
    .A2(_03153_),
    .B1(_03460_),
    .B2(_03461_),
    .X(cpu_rdata[56]));
 sky130_fd_sc_hd__o21a_2 _06002_ (.A1(\data_array.rdata0[57] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03462_));
 sky130_fd_sc_hd__a21o_2 _06003_ (.A1(\data_array.rdata1[57] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03463_));
 sky130_fd_sc_hd__a22o_2 _06004_ (.A1(mem_rdata[57]),
    .A2(_03153_),
    .B1(_03462_),
    .B2(_03463_),
    .X(cpu_rdata[57]));
 sky130_fd_sc_hd__o21a_2 _06005_ (.A1(\data_array.rdata0[58] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03464_));
 sky130_fd_sc_hd__a21o_2 _06006_ (.A1(\data_array.rdata1[58] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03465_));
 sky130_fd_sc_hd__a22o_2 _06007_ (.A1(mem_rdata[58]),
    .A2(_03153_),
    .B1(_03464_),
    .B2(_03465_),
    .X(cpu_rdata[58]));
 sky130_fd_sc_hd__o21a_2 _06008_ (.A1(\data_array.rdata0[59] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03466_));
 sky130_fd_sc_hd__a21o_2 _06009_ (.A1(\data_array.rdata1[59] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03467_));
 sky130_fd_sc_hd__a22o_2 _06010_ (.A1(mem_rdata[59]),
    .A2(_03153_),
    .B1(_03466_),
    .B2(_03467_),
    .X(cpu_rdata[59]));
 sky130_fd_sc_hd__o21a_2 _06011_ (.A1(\data_array.rdata0[60] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03468_));
 sky130_fd_sc_hd__a21o_2 _06012_ (.A1(\data_array.rdata1[60] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03469_));
 sky130_fd_sc_hd__a22o_2 _06013_ (.A1(mem_rdata[60]),
    .A2(_03153_),
    .B1(_03468_),
    .B2(_03469_),
    .X(cpu_rdata[60]));
 sky130_fd_sc_hd__o21a_2 _06014_ (.A1(\data_array.rdata0[61] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03470_));
 sky130_fd_sc_hd__a21o_2 _06015_ (.A1(\data_array.rdata1[61] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03471_));
 sky130_fd_sc_hd__a22o_2 _06016_ (.A1(mem_rdata[61]),
    .A2(_03153_),
    .B1(_03470_),
    .B2(_03471_),
    .X(cpu_rdata[61]));
 sky130_fd_sc_hd__o21a_2 _06017_ (.A1(\data_array.rdata0[62] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03472_));
 sky130_fd_sc_hd__a21o_2 _06018_ (.A1(\data_array.rdata1[62] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03473_));
 sky130_fd_sc_hd__a22o_2 _06019_ (.A1(mem_rdata[62]),
    .A2(_03153_),
    .B1(_03472_),
    .B2(_03473_),
    .X(cpu_rdata[62]));
 sky130_fd_sc_hd__o21a_2 _06020_ (.A1(\data_array.rdata0[63] ),
    .A2(_03213_),
    .B1(_03154_),
    .X(_03474_));
 sky130_fd_sc_hd__a21o_2 _06021_ (.A1(\data_array.rdata1[63] ),
    .A2(_03315_),
    .B1(_03236_),
    .X(_03475_));
 sky130_fd_sc_hd__a22o_2 _06022_ (.A1(mem_rdata[63]),
    .A2(_03153_),
    .B1(_03474_),
    .B2(_03475_),
    .X(cpu_rdata[63]));
 sky130_fd_sc_hd__and2_2 _06023_ (.A(mem_read),
    .B(cpu_addr[0]),
    .X(mem_addr[0]));
 sky130_fd_sc_hd__and2_2 _06024_ (.A(mem_read),
    .B(cpu_addr[1]),
    .X(mem_addr[1]));
 sky130_fd_sc_hd__and2_2 _06025_ (.A(mem_read),
    .B(cpu_addr[2]),
    .X(mem_addr[2]));
 sky130_fd_sc_hd__and2b_2 _06026_ (.A_N(\fsm.lru_out ),
    .B(mem_write),
    .X(_03476_));
 sky130_fd_sc_hd__and3b_2 _06027_ (.A_N(\fsm.lru_out ),
    .B(\fsm.state[5] ),
    .C(\fsm.valid0 ),
    .X(_03477_));
 sky130_fd_sc_hd__or2_2 _06028_ (.A(_03476_),
    .B(_03477_),
    .X(_03478_));
 sky130_fd_sc_hd__and3_2 _06029_ (.A(\fsm.lru_out ),
    .B(\fsm.valid1 ),
    .C(\fsm.state[5] ),
    .X(_03479_));
 sky130_fd_sc_hd__or2_2 _06030_ (.A(_03476_),
    .B(_03479_),
    .X(_03480_));
 sky130_fd_sc_hd__o31a_2 _06031_ (.A1(mem_read),
    .A2(_03477_),
    .A3(_03480_),
    .B1(cpu_addr[3]),
    .X(mem_addr[3]));
 sky130_fd_sc_hd__o31a_2 _06032_ (.A1(mem_read),
    .A2(_03477_),
    .A3(_03480_),
    .B1(cpu_addr[4]),
    .X(mem_addr[4]));
 sky130_fd_sc_hd__o31a_2 _06033_ (.A1(mem_read),
    .A2(_03477_),
    .A3(_03480_),
    .B1(cpu_addr[5]),
    .X(mem_addr[5]));
 sky130_fd_sc_hd__o31a_2 _06034_ (.A1(mem_read),
    .A2(_03477_),
    .A3(_03480_),
    .B1(cpu_addr[6]),
    .X(mem_addr[6]));
 sky130_fd_sc_hd__a22o_2 _06035_ (.A1(mem_read),
    .A2(cpu_addr[7]),
    .B1(\fsm.tag_out1[0] ),
    .B2(_03479_),
    .X(_03481_));
 sky130_fd_sc_hd__a21o_2 _06036_ (.A1(\fsm.tag_out0[0] ),
    .A2(_03478_),
    .B1(_03481_),
    .X(mem_addr[7]));
 sky130_fd_sc_hd__a22o_2 _06037_ (.A1(mem_read),
    .A2(cpu_addr[8]),
    .B1(\fsm.tag_out1[1] ),
    .B2(_03479_),
    .X(_03482_));
 sky130_fd_sc_hd__a21o_2 _06038_ (.A1(\fsm.tag_out0[1] ),
    .A2(_03478_),
    .B1(_03482_),
    .X(mem_addr[8]));
 sky130_fd_sc_hd__a22o_2 _06039_ (.A1(mem_read),
    .A2(cpu_addr[9]),
    .B1(\fsm.tag_out1[2] ),
    .B2(_03479_),
    .X(_03483_));
 sky130_fd_sc_hd__a21o_2 _06040_ (.A1(\fsm.tag_out0[2] ),
    .A2(_03478_),
    .B1(_03483_),
    .X(mem_addr[9]));
 sky130_fd_sc_hd__a22o_2 _06041_ (.A1(mem_read),
    .A2(cpu_addr[10]),
    .B1(\fsm.tag_out1[3] ),
    .B2(_03479_),
    .X(_03484_));
 sky130_fd_sc_hd__a21o_2 _06042_ (.A1(\fsm.tag_out0[3] ),
    .A2(_03478_),
    .B1(_03484_),
    .X(mem_addr[10]));
 sky130_fd_sc_hd__a22o_2 _06043_ (.A1(mem_read),
    .A2(cpu_addr[11]),
    .B1(\fsm.tag_out1[4] ),
    .B2(_03479_),
    .X(_03485_));
 sky130_fd_sc_hd__a21o_2 _06044_ (.A1(\fsm.tag_out0[4] ),
    .A2(_03478_),
    .B1(_03485_),
    .X(mem_addr[11]));
 sky130_fd_sc_hd__a22o_2 _06045_ (.A1(mem_read),
    .A2(cpu_addr[12]),
    .B1(\fsm.tag_out1[5] ),
    .B2(_03479_),
    .X(_03486_));
 sky130_fd_sc_hd__a21o_2 _06046_ (.A1(\fsm.tag_out0[5] ),
    .A2(_03478_),
    .B1(_03486_),
    .X(mem_addr[12]));
 sky130_fd_sc_hd__a22o_2 _06047_ (.A1(mem_read),
    .A2(cpu_addr[13]),
    .B1(\fsm.tag_out1[6] ),
    .B2(_03479_),
    .X(_03487_));
 sky130_fd_sc_hd__a21o_2 _06048_ (.A1(\fsm.tag_out0[6] ),
    .A2(_03478_),
    .B1(_03487_),
    .X(mem_addr[13]));
 sky130_fd_sc_hd__a22o_2 _06049_ (.A1(mem_read),
    .A2(cpu_addr[14]),
    .B1(\fsm.tag_out1[7] ),
    .B2(_03479_),
    .X(_03488_));
 sky130_fd_sc_hd__a21o_2 _06050_ (.A1(\fsm.tag_out0[7] ),
    .A2(_03478_),
    .B1(_03488_),
    .X(mem_addr[14]));
 sky130_fd_sc_hd__a22o_2 _06051_ (.A1(mem_read),
    .A2(cpu_addr[15]),
    .B1(\fsm.tag_out1[8] ),
    .B2(_03479_),
    .X(_03489_));
 sky130_fd_sc_hd__a21o_2 _06052_ (.A1(\fsm.tag_out0[8] ),
    .A2(_03478_),
    .B1(_03489_),
    .X(mem_addr[15]));
 sky130_fd_sc_hd__a22o_2 _06053_ (.A1(mem_read),
    .A2(cpu_addr[16]),
    .B1(\fsm.tag_out1[9] ),
    .B2(_03479_),
    .X(_03490_));
 sky130_fd_sc_hd__a21o_2 _06054_ (.A1(\fsm.tag_out0[9] ),
    .A2(_03478_),
    .B1(_03490_),
    .X(mem_addr[16]));
 sky130_fd_sc_hd__a22o_2 _06055_ (.A1(mem_read),
    .A2(cpu_addr[17]),
    .B1(\fsm.tag_out1[10] ),
    .B2(_03479_),
    .X(_03491_));
 sky130_fd_sc_hd__a21o_2 _06056_ (.A1(\fsm.tag_out0[10] ),
    .A2(_03478_),
    .B1(_03491_),
    .X(mem_addr[17]));
 sky130_fd_sc_hd__a22o_2 _06057_ (.A1(mem_read),
    .A2(cpu_addr[18]),
    .B1(\fsm.tag_out1[11] ),
    .B2(_03479_),
    .X(_03492_));
 sky130_fd_sc_hd__a21o_2 _06058_ (.A1(\fsm.tag_out0[11] ),
    .A2(_03478_),
    .B1(_03492_),
    .X(mem_addr[18]));
 sky130_fd_sc_hd__a22o_2 _06059_ (.A1(mem_read),
    .A2(cpu_addr[19]),
    .B1(\fsm.tag_out1[12] ),
    .B2(_03479_),
    .X(_03493_));
 sky130_fd_sc_hd__a21o_2 _06060_ (.A1(\fsm.tag_out0[12] ),
    .A2(_03478_),
    .B1(_03493_),
    .X(mem_addr[19]));
 sky130_fd_sc_hd__a22o_2 _06061_ (.A1(mem_read),
    .A2(cpu_addr[20]),
    .B1(\fsm.tag_out1[13] ),
    .B2(_03479_),
    .X(_03494_));
 sky130_fd_sc_hd__a21o_2 _06062_ (.A1(\fsm.tag_out0[13] ),
    .A2(_03478_),
    .B1(_03494_),
    .X(mem_addr[20]));
 sky130_fd_sc_hd__a22o_2 _06063_ (.A1(mem_read),
    .A2(cpu_addr[21]),
    .B1(\fsm.tag_out1[14] ),
    .B2(_03479_),
    .X(_03495_));
 sky130_fd_sc_hd__a21o_2 _06064_ (.A1(\fsm.tag_out0[14] ),
    .A2(_03478_),
    .B1(_03495_),
    .X(mem_addr[21]));
 sky130_fd_sc_hd__a22o_2 _06065_ (.A1(mem_read),
    .A2(cpu_addr[22]),
    .B1(\fsm.tag_out1[15] ),
    .B2(_03479_),
    .X(_03496_));
 sky130_fd_sc_hd__a21o_2 _06066_ (.A1(\fsm.tag_out0[15] ),
    .A2(_03478_),
    .B1(_03496_),
    .X(mem_addr[22]));
 sky130_fd_sc_hd__a22o_2 _06067_ (.A1(mem_read),
    .A2(cpu_addr[23]),
    .B1(\fsm.tag_out1[16] ),
    .B2(_03479_),
    .X(_03497_));
 sky130_fd_sc_hd__a21o_2 _06068_ (.A1(\fsm.tag_out0[16] ),
    .A2(_03478_),
    .B1(_03497_),
    .X(mem_addr[23]));
 sky130_fd_sc_hd__a22o_2 _06069_ (.A1(mem_read),
    .A2(cpu_addr[24]),
    .B1(\fsm.tag_out1[17] ),
    .B2(_03479_),
    .X(_03498_));
 sky130_fd_sc_hd__a21o_2 _06070_ (.A1(\fsm.tag_out0[17] ),
    .A2(_03478_),
    .B1(_03498_),
    .X(mem_addr[24]));
 sky130_fd_sc_hd__a22o_2 _06071_ (.A1(mem_read),
    .A2(cpu_addr[25]),
    .B1(\fsm.tag_out1[18] ),
    .B2(_03479_),
    .X(_03499_));
 sky130_fd_sc_hd__a21o_2 _06072_ (.A1(\fsm.tag_out0[18] ),
    .A2(_03478_),
    .B1(_03499_),
    .X(mem_addr[25]));
 sky130_fd_sc_hd__a22o_2 _06073_ (.A1(mem_read),
    .A2(cpu_addr[26]),
    .B1(\fsm.tag_out1[19] ),
    .B2(_03479_),
    .X(_03500_));
 sky130_fd_sc_hd__a21o_2 _06074_ (.A1(\fsm.tag_out0[19] ),
    .A2(_03478_),
    .B1(_03500_),
    .X(mem_addr[26]));
 sky130_fd_sc_hd__a22o_2 _06075_ (.A1(mem_read),
    .A2(cpu_addr[27]),
    .B1(\fsm.tag_out1[20] ),
    .B2(_03479_),
    .X(_03501_));
 sky130_fd_sc_hd__a21o_2 _06076_ (.A1(\fsm.tag_out0[20] ),
    .A2(_03478_),
    .B1(_03501_),
    .X(mem_addr[27]));
 sky130_fd_sc_hd__a22o_2 _06077_ (.A1(mem_read),
    .A2(cpu_addr[28]),
    .B1(\fsm.tag_out1[21] ),
    .B2(_03479_),
    .X(_03502_));
 sky130_fd_sc_hd__a21o_2 _06078_ (.A1(\fsm.tag_out0[21] ),
    .A2(_03478_),
    .B1(_03502_),
    .X(mem_addr[28]));
 sky130_fd_sc_hd__a22o_2 _06079_ (.A1(mem_read),
    .A2(cpu_addr[29]),
    .B1(\fsm.tag_out1[22] ),
    .B2(_03479_),
    .X(_03503_));
 sky130_fd_sc_hd__a21o_2 _06080_ (.A1(\fsm.tag_out0[22] ),
    .A2(_03478_),
    .B1(_03503_),
    .X(mem_addr[29]));
 sky130_fd_sc_hd__a22o_2 _06081_ (.A1(mem_read),
    .A2(cpu_addr[30]),
    .B1(\fsm.tag_out1[23] ),
    .B2(_03479_),
    .X(_03504_));
 sky130_fd_sc_hd__a21o_2 _06082_ (.A1(\fsm.tag_out0[23] ),
    .A2(_03478_),
    .B1(_03504_),
    .X(mem_addr[30]));
 sky130_fd_sc_hd__a22o_2 _06083_ (.A1(mem_read),
    .A2(cpu_addr[31]),
    .B1(\fsm.tag_out1[24] ),
    .B2(_03479_),
    .X(_03505_));
 sky130_fd_sc_hd__a21o_2 _06084_ (.A1(\fsm.tag_out0[24] ),
    .A2(_03478_),
    .B1(_03505_),
    .X(mem_addr[31]));
 sky130_fd_sc_hd__a22o_2 _06085_ (.A1(\data_array.rdata0[0] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[0] ),
    .X(mem_wdata[0]));
 sky130_fd_sc_hd__a22o_2 _06086_ (.A1(\data_array.rdata0[1] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[1] ),
    .X(mem_wdata[1]));
 sky130_fd_sc_hd__a22o_2 _06087_ (.A1(\data_array.rdata0[2] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[2] ),
    .X(mem_wdata[2]));
 sky130_fd_sc_hd__a22o_2 _06088_ (.A1(\data_array.rdata0[3] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[3] ),
    .X(mem_wdata[3]));
 sky130_fd_sc_hd__a22o_2 _06089_ (.A1(\data_array.rdata0[4] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[4] ),
    .X(mem_wdata[4]));
 sky130_fd_sc_hd__a22o_2 _06090_ (.A1(\data_array.rdata0[5] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[5] ),
    .X(mem_wdata[5]));
 sky130_fd_sc_hd__a22o_2 _06091_ (.A1(\data_array.rdata0[6] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[6] ),
    .X(mem_wdata[6]));
 sky130_fd_sc_hd__a22o_2 _06092_ (.A1(\data_array.rdata0[7] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[7] ),
    .X(mem_wdata[7]));
 sky130_fd_sc_hd__a22o_2 _06093_ (.A1(\data_array.rdata0[8] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[8] ),
    .X(mem_wdata[8]));
 sky130_fd_sc_hd__a22o_2 _06094_ (.A1(\data_array.rdata0[9] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[9] ),
    .X(mem_wdata[9]));
 sky130_fd_sc_hd__a22o_2 _06095_ (.A1(\data_array.rdata0[10] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[10] ),
    .X(mem_wdata[10]));
 sky130_fd_sc_hd__a22o_2 _06096_ (.A1(\data_array.rdata0[11] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[11] ),
    .X(mem_wdata[11]));
 sky130_fd_sc_hd__a22o_2 _06097_ (.A1(\data_array.rdata0[12] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[12] ),
    .X(mem_wdata[12]));
 sky130_fd_sc_hd__a22o_2 _06098_ (.A1(\data_array.rdata0[13] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[13] ),
    .X(mem_wdata[13]));
 sky130_fd_sc_hd__a22o_2 _06099_ (.A1(\data_array.rdata0[14] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[14] ),
    .X(mem_wdata[14]));
 sky130_fd_sc_hd__a22o_2 _06100_ (.A1(\data_array.rdata0[15] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[15] ),
    .X(mem_wdata[15]));
 sky130_fd_sc_hd__a22o_2 _06101_ (.A1(\data_array.rdata0[16] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[16] ),
    .X(mem_wdata[16]));
 sky130_fd_sc_hd__a22o_2 _06102_ (.A1(\data_array.rdata0[17] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[17] ),
    .X(mem_wdata[17]));
 sky130_fd_sc_hd__a22o_2 _06103_ (.A1(\data_array.rdata0[18] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[18] ),
    .X(mem_wdata[18]));
 sky130_fd_sc_hd__a22o_2 _06104_ (.A1(\data_array.rdata0[19] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[19] ),
    .X(mem_wdata[19]));
 sky130_fd_sc_hd__a22o_2 _06105_ (.A1(\data_array.rdata0[20] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[20] ),
    .X(mem_wdata[20]));
 sky130_fd_sc_hd__a22o_2 _06106_ (.A1(\data_array.rdata0[21] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[21] ),
    .X(mem_wdata[21]));
 sky130_fd_sc_hd__a22o_2 _06107_ (.A1(\data_array.rdata0[22] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[22] ),
    .X(mem_wdata[22]));
 sky130_fd_sc_hd__a22o_2 _06108_ (.A1(\data_array.rdata0[23] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[23] ),
    .X(mem_wdata[23]));
 sky130_fd_sc_hd__a22o_2 _06109_ (.A1(\data_array.rdata0[24] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[24] ),
    .X(mem_wdata[24]));
 sky130_fd_sc_hd__a22o_2 _06110_ (.A1(\data_array.rdata0[25] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[25] ),
    .X(mem_wdata[25]));
 sky130_fd_sc_hd__a22o_2 _06111_ (.A1(\data_array.rdata0[26] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[26] ),
    .X(mem_wdata[26]));
 sky130_fd_sc_hd__a22o_2 _06112_ (.A1(\data_array.rdata0[27] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[27] ),
    .X(mem_wdata[27]));
 sky130_fd_sc_hd__a22o_2 _06113_ (.A1(\data_array.rdata0[28] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[28] ),
    .X(mem_wdata[28]));
 sky130_fd_sc_hd__a22o_2 _06114_ (.A1(\data_array.rdata0[29] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[29] ),
    .X(mem_wdata[29]));
 sky130_fd_sc_hd__a22o_2 _06115_ (.A1(\data_array.rdata0[30] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[30] ),
    .X(mem_wdata[30]));
 sky130_fd_sc_hd__a22o_2 _06116_ (.A1(\data_array.rdata0[31] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[31] ),
    .X(mem_wdata[31]));
 sky130_fd_sc_hd__a22o_2 _06117_ (.A1(\data_array.rdata0[32] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[32] ),
    .X(mem_wdata[32]));
 sky130_fd_sc_hd__a22o_2 _06118_ (.A1(\data_array.rdata0[33] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[33] ),
    .X(mem_wdata[33]));
 sky130_fd_sc_hd__a22o_2 _06119_ (.A1(\data_array.rdata0[34] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[34] ),
    .X(mem_wdata[34]));
 sky130_fd_sc_hd__a22o_2 _06120_ (.A1(\data_array.rdata0[35] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[35] ),
    .X(mem_wdata[35]));
 sky130_fd_sc_hd__a22o_2 _06121_ (.A1(\data_array.rdata0[36] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[36] ),
    .X(mem_wdata[36]));
 sky130_fd_sc_hd__a22o_2 _06122_ (.A1(\data_array.rdata0[37] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[37] ),
    .X(mem_wdata[37]));
 sky130_fd_sc_hd__a22o_2 _06123_ (.A1(\data_array.rdata0[38] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[38] ),
    .X(mem_wdata[38]));
 sky130_fd_sc_hd__a22o_2 _06124_ (.A1(\data_array.rdata0[39] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[39] ),
    .X(mem_wdata[39]));
 sky130_fd_sc_hd__a22o_2 _06125_ (.A1(\data_array.rdata0[40] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[40] ),
    .X(mem_wdata[40]));
 sky130_fd_sc_hd__a22o_2 _06126_ (.A1(\data_array.rdata0[41] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[41] ),
    .X(mem_wdata[41]));
 sky130_fd_sc_hd__a22o_2 _06127_ (.A1(\data_array.rdata0[42] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[42] ),
    .X(mem_wdata[42]));
 sky130_fd_sc_hd__a22o_2 _06128_ (.A1(\data_array.rdata0[43] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[43] ),
    .X(mem_wdata[43]));
 sky130_fd_sc_hd__a22o_2 _06129_ (.A1(\data_array.rdata0[44] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[44] ),
    .X(mem_wdata[44]));
 sky130_fd_sc_hd__a22o_2 _06130_ (.A1(\data_array.rdata0[45] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[45] ),
    .X(mem_wdata[45]));
 sky130_fd_sc_hd__a22o_2 _06131_ (.A1(\data_array.rdata0[46] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[46] ),
    .X(mem_wdata[46]));
 sky130_fd_sc_hd__a22o_2 _06132_ (.A1(\data_array.rdata0[47] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[47] ),
    .X(mem_wdata[47]));
 sky130_fd_sc_hd__a22o_2 _06133_ (.A1(\data_array.rdata0[48] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[48] ),
    .X(mem_wdata[48]));
 sky130_fd_sc_hd__a22o_2 _06134_ (.A1(\data_array.rdata0[49] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[49] ),
    .X(mem_wdata[49]));
 sky130_fd_sc_hd__a22o_2 _06135_ (.A1(\data_array.rdata0[50] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[50] ),
    .X(mem_wdata[50]));
 sky130_fd_sc_hd__a22o_2 _06136_ (.A1(\data_array.rdata0[51] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[51] ),
    .X(mem_wdata[51]));
 sky130_fd_sc_hd__a22o_2 _06137_ (.A1(\data_array.rdata0[52] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[52] ),
    .X(mem_wdata[52]));
 sky130_fd_sc_hd__a22o_2 _06138_ (.A1(\data_array.rdata0[53] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[53] ),
    .X(mem_wdata[53]));
 sky130_fd_sc_hd__a22o_2 _06139_ (.A1(\data_array.rdata0[54] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[54] ),
    .X(mem_wdata[54]));
 sky130_fd_sc_hd__a22o_2 _06140_ (.A1(\data_array.rdata0[55] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[55] ),
    .X(mem_wdata[55]));
 sky130_fd_sc_hd__a22o_2 _06141_ (.A1(\data_array.rdata0[56] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[56] ),
    .X(mem_wdata[56]));
 sky130_fd_sc_hd__a22o_2 _06142_ (.A1(\data_array.rdata0[57] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[57] ),
    .X(mem_wdata[57]));
 sky130_fd_sc_hd__a22o_2 _06143_ (.A1(\data_array.rdata0[58] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[58] ),
    .X(mem_wdata[58]));
 sky130_fd_sc_hd__a22o_2 _06144_ (.A1(\data_array.rdata0[59] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[59] ),
    .X(mem_wdata[59]));
 sky130_fd_sc_hd__a22o_2 _06145_ (.A1(\data_array.rdata0[60] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[60] ),
    .X(mem_wdata[60]));
 sky130_fd_sc_hd__a22o_2 _06146_ (.A1(\data_array.rdata0[61] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[61] ),
    .X(mem_wdata[61]));
 sky130_fd_sc_hd__a22o_2 _06147_ (.A1(\data_array.rdata0[62] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[62] ),
    .X(mem_wdata[62]));
 sky130_fd_sc_hd__a22o_2 _06148_ (.A1(\data_array.rdata0[63] ),
    .A2(_03477_),
    .B1(_03480_),
    .B2(\data_array.rdata1[63] ),
    .X(mem_wdata[63]));
 sky130_fd_sc_hd__and2b_2 _06149_ (.A_N(cpu_addr[5]),
    .B(cpu_addr[6]),
    .X(_03506_));
 sky130_fd_sc_hd__nand2b_2 _06150_ (.A_N(cpu_addr[5]),
    .B(cpu_addr[6]),
    .Y(_03507_));
 sky130_fd_sc_hd__and2b_2 _06151_ (.A_N(cpu_addr[4]),
    .B(cpu_addr[3]),
    .X(_03508_));
 sky130_fd_sc_hd__nand2b_2 _06152_ (.A_N(cpu_addr[4]),
    .B(cpu_addr[3]),
    .Y(_03509_));
 sky130_fd_sc_hd__and2b_2 _06153_ (.A_N(cpu_addr[3]),
    .B(cpu_addr[4]),
    .X(_03510_));
 sky130_fd_sc_hd__nand2b_2 _06154_ (.A_N(cpu_addr[3]),
    .B(cpu_addr[4]),
    .Y(_03511_));
 sky130_fd_sc_hd__a22o_2 _06155_ (.A1(\tag_array.valid0[9] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.valid0[10] ),
    .X(_03512_));
 sky130_fd_sc_hd__nor2_2 _06156_ (.A(cpu_addr[3]),
    .B(cpu_addr[4]),
    .Y(_03513_));
 sky130_fd_sc_hd__or2_2 _06157_ (.A(cpu_addr[3]),
    .B(cpu_addr[4]),
    .X(_03514_));
 sky130_fd_sc_hd__and2_2 _06158_ (.A(cpu_addr[3]),
    .B(cpu_addr[4]),
    .X(_03515_));
 sky130_fd_sc_hd__nand2_2 _06159_ (.A(cpu_addr[3]),
    .B(cpu_addr[4]),
    .Y(_03516_));
 sky130_fd_sc_hd__a221o_2 _06160_ (.A1(\tag_array.valid0[8] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.valid0[11] ),
    .C1(_03512_),
    .X(_03517_));
 sky130_fd_sc_hd__nor2_2 _06161_ (.A(cpu_addr[5]),
    .B(cpu_addr[6]),
    .Y(_03518_));
 sky130_fd_sc_hd__or2_2 _06162_ (.A(cpu_addr[5]),
    .B(cpu_addr[6]),
    .X(_03519_));
 sky130_fd_sc_hd__a22o_2 _06163_ (.A1(\tag_array.valid0[1] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.valid0[2] ),
    .X(_03520_));
 sky130_fd_sc_hd__a221o_2 _06164_ (.A1(\tag_array.valid0[0] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.valid0[3] ),
    .C1(_03520_),
    .X(_03521_));
 sky130_fd_sc_hd__and2_2 _06165_ (.A(cpu_addr[5]),
    .B(cpu_addr[6]),
    .X(_03522_));
 sky130_fd_sc_hd__nand2_2 _06166_ (.A(cpu_addr[5]),
    .B(cpu_addr[6]),
    .Y(_03523_));
 sky130_fd_sc_hd__a22o_2 _06167_ (.A1(\tag_array.valid0[13] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.valid0[14] ),
    .X(_03524_));
 sky130_fd_sc_hd__a221o_2 _06168_ (.A1(\tag_array.valid0[12] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.valid0[15] ),
    .C1(_03524_),
    .X(_03525_));
 sky130_fd_sc_hd__and2b_2 _06169_ (.A_N(cpu_addr[6]),
    .B(cpu_addr[5]),
    .X(_03526_));
 sky130_fd_sc_hd__nand2b_2 _06170_ (.A_N(cpu_addr[6]),
    .B(cpu_addr[5]),
    .Y(_03527_));
 sky130_fd_sc_hd__a22o_2 _06171_ (.A1(\tag_array.valid0[5] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.valid0[6] ),
    .X(_03528_));
 sky130_fd_sc_hd__a221o_2 _06172_ (.A1(\tag_array.valid0[4] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.valid0[7] ),
    .C1(_03528_),
    .X(_03529_));
 sky130_fd_sc_hd__a22o_2 _06173_ (.A1(_03506_),
    .A2(_03517_),
    .B1(_03522_),
    .B2(_03525_),
    .X(_03530_));
 sky130_fd_sc_hd__a22o_2 _06174_ (.A1(_03518_),
    .A2(_03521_),
    .B1(_03526_),
    .B2(_03529_),
    .X(_03531_));
 sky130_fd_sc_hd__or2_2 _06175_ (.A(_03530_),
    .B(_03531_),
    .X(_00181_));
 sky130_fd_sc_hd__a22o_2 _06176_ (.A1(\tag_array.valid1[13] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.valid1[14] ),
    .X(_03532_));
 sky130_fd_sc_hd__a221o_2 _06177_ (.A1(\tag_array.valid1[12] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.valid1[15] ),
    .C1(_03532_),
    .X(_03533_));
 sky130_fd_sc_hd__a22o_2 _06178_ (.A1(\tag_array.valid1[1] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.valid1[2] ),
    .X(_03534_));
 sky130_fd_sc_hd__a221o_2 _06179_ (.A1(\tag_array.valid1[0] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.valid1[3] ),
    .C1(_03534_),
    .X(_03535_));
 sky130_fd_sc_hd__a22o_2 _06180_ (.A1(\tag_array.valid1[9] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.valid1[10] ),
    .X(_03536_));
 sky130_fd_sc_hd__a221o_2 _06181_ (.A1(\tag_array.valid1[8] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.valid1[11] ),
    .C1(_03536_),
    .X(_03537_));
 sky130_fd_sc_hd__a22o_2 _06182_ (.A1(\tag_array.valid1[5] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.valid1[6] ),
    .X(_03538_));
 sky130_fd_sc_hd__a221o_2 _06183_ (.A1(\tag_array.valid1[4] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.valid1[7] ),
    .C1(_03538_),
    .X(_03539_));
 sky130_fd_sc_hd__a22o_2 _06184_ (.A1(_03522_),
    .A2(_03533_),
    .B1(_03537_),
    .B2(_03506_),
    .X(_03540_));
 sky130_fd_sc_hd__a22o_2 _06185_ (.A1(_03518_),
    .A2(_03535_),
    .B1(_03539_),
    .B2(_03526_),
    .X(_03541_));
 sky130_fd_sc_hd__or2_2 _06186_ (.A(_03540_),
    .B(_03541_),
    .X(_00182_));
 sky130_fd_sc_hd__a22o_2 _06187_ (.A1(\tag_array.tag0[9][0] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[10][0] ),
    .X(_03542_));
 sky130_fd_sc_hd__a221o_2 _06188_ (.A1(\tag_array.tag0[8][0] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[11][0] ),
    .C1(_03542_),
    .X(_03543_));
 sky130_fd_sc_hd__a22o_2 _06189_ (.A1(\tag_array.tag0[5][0] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[6][0] ),
    .X(_03544_));
 sky130_fd_sc_hd__a221o_2 _06190_ (.A1(\tag_array.tag0[4][0] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[7][0] ),
    .C1(_03544_),
    .X(_03545_));
 sky130_fd_sc_hd__a22o_2 _06191_ (.A1(\tag_array.tag0[13][0] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[14][0] ),
    .X(_03546_));
 sky130_fd_sc_hd__a221o_2 _06192_ (.A1(\tag_array.tag0[12][0] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[15][0] ),
    .C1(_03546_),
    .X(_03547_));
 sky130_fd_sc_hd__a22o_2 _06193_ (.A1(\tag_array.tag0[1][0] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[2][0] ),
    .X(_03548_));
 sky130_fd_sc_hd__a221o_2 _06194_ (.A1(\tag_array.tag0[0][0] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[3][0] ),
    .C1(_03548_),
    .X(_03549_));
 sky130_fd_sc_hd__a22o_2 _06195_ (.A1(_03506_),
    .A2(_03543_),
    .B1(_03547_),
    .B2(_03522_),
    .X(_03550_));
 sky130_fd_sc_hd__a22o_2 _06196_ (.A1(_03526_),
    .A2(_03545_),
    .B1(_03549_),
    .B2(_03518_),
    .X(_03551_));
 sky130_fd_sc_hd__or2_2 _06197_ (.A(_03550_),
    .B(_03551_),
    .X(_00131_));
 sky130_fd_sc_hd__a22o_2 _06198_ (.A1(\tag_array.tag0[9][1] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[10][1] ),
    .X(_03552_));
 sky130_fd_sc_hd__a221o_2 _06199_ (.A1(\tag_array.tag0[8][1] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[11][1] ),
    .C1(_03552_),
    .X(_03553_));
 sky130_fd_sc_hd__a22o_2 _06200_ (.A1(\tag_array.tag0[5][1] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[6][1] ),
    .X(_03554_));
 sky130_fd_sc_hd__a221o_2 _06201_ (.A1(\tag_array.tag0[4][1] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[7][1] ),
    .C1(_03554_),
    .X(_03555_));
 sky130_fd_sc_hd__a22o_2 _06202_ (.A1(\tag_array.tag0[13][1] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[14][1] ),
    .X(_03556_));
 sky130_fd_sc_hd__a221o_2 _06203_ (.A1(\tag_array.tag0[12][1] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[15][1] ),
    .C1(_03556_),
    .X(_03557_));
 sky130_fd_sc_hd__a22o_2 _06204_ (.A1(\tag_array.tag0[1][1] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[2][1] ),
    .X(_03558_));
 sky130_fd_sc_hd__a221o_2 _06205_ (.A1(\tag_array.tag0[0][1] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[3][1] ),
    .C1(_03558_),
    .X(_03559_));
 sky130_fd_sc_hd__a22o_2 _06206_ (.A1(_03506_),
    .A2(_03553_),
    .B1(_03557_),
    .B2(_03522_),
    .X(_03560_));
 sky130_fd_sc_hd__a22o_2 _06207_ (.A1(_03526_),
    .A2(_03555_),
    .B1(_03559_),
    .B2(_03518_),
    .X(_03561_));
 sky130_fd_sc_hd__or2_2 _06208_ (.A(_03560_),
    .B(_03561_),
    .X(_00142_));
 sky130_fd_sc_hd__a22o_2 _06209_ (.A1(\tag_array.tag0[9][2] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[10][2] ),
    .X(_03562_));
 sky130_fd_sc_hd__a221o_2 _06210_ (.A1(\tag_array.tag0[8][2] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[11][2] ),
    .C1(_03562_),
    .X(_03563_));
 sky130_fd_sc_hd__a22o_2 _06211_ (.A1(\tag_array.tag0[5][2] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[6][2] ),
    .X(_03564_));
 sky130_fd_sc_hd__a221o_2 _06212_ (.A1(\tag_array.tag0[4][2] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[7][2] ),
    .C1(_03564_),
    .X(_03565_));
 sky130_fd_sc_hd__a22o_2 _06213_ (.A1(\tag_array.tag0[13][2] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[14][2] ),
    .X(_03566_));
 sky130_fd_sc_hd__a221o_2 _06214_ (.A1(\tag_array.tag0[12][2] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[15][2] ),
    .C1(_03566_),
    .X(_03567_));
 sky130_fd_sc_hd__a22o_2 _06215_ (.A1(\tag_array.tag0[1][2] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[2][2] ),
    .X(_03568_));
 sky130_fd_sc_hd__a221o_2 _06216_ (.A1(\tag_array.tag0[0][2] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[3][2] ),
    .C1(_03568_),
    .X(_03569_));
 sky130_fd_sc_hd__a22o_2 _06217_ (.A1(_03506_),
    .A2(_03563_),
    .B1(_03567_),
    .B2(_03522_),
    .X(_03570_));
 sky130_fd_sc_hd__a22o_2 _06218_ (.A1(_03526_),
    .A2(_03565_),
    .B1(_03569_),
    .B2(_03518_),
    .X(_03571_));
 sky130_fd_sc_hd__or2_2 _06219_ (.A(_03570_),
    .B(_03571_),
    .X(_00148_));
 sky130_fd_sc_hd__a22o_2 _06220_ (.A1(\tag_array.tag0[13][3] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[14][3] ),
    .X(_03572_));
 sky130_fd_sc_hd__a221o_2 _06221_ (.A1(\tag_array.tag0[12][3] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[15][3] ),
    .C1(_03572_),
    .X(_03573_));
 sky130_fd_sc_hd__a22o_2 _06222_ (.A1(\tag_array.tag0[1][3] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[2][3] ),
    .X(_03574_));
 sky130_fd_sc_hd__a221o_2 _06223_ (.A1(\tag_array.tag0[0][3] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[3][3] ),
    .C1(_03574_),
    .X(_03575_));
 sky130_fd_sc_hd__a22o_2 _06224_ (.A1(\tag_array.tag0[9][3] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[10][3] ),
    .X(_03576_));
 sky130_fd_sc_hd__a221o_2 _06225_ (.A1(\tag_array.tag0[8][3] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[11][3] ),
    .C1(_03576_),
    .X(_03577_));
 sky130_fd_sc_hd__a22o_2 _06226_ (.A1(\tag_array.tag0[5][3] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[6][3] ),
    .X(_03578_));
 sky130_fd_sc_hd__a221o_2 _06227_ (.A1(\tag_array.tag0[4][3] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[7][3] ),
    .C1(_03578_),
    .X(_03579_));
 sky130_fd_sc_hd__a22o_2 _06228_ (.A1(_03522_),
    .A2(_03573_),
    .B1(_03577_),
    .B2(_03506_),
    .X(_03580_));
 sky130_fd_sc_hd__a22o_2 _06229_ (.A1(_03518_),
    .A2(_03575_),
    .B1(_03579_),
    .B2(_03526_),
    .X(_03581_));
 sky130_fd_sc_hd__or2_2 _06230_ (.A(_03580_),
    .B(_03581_),
    .X(_00149_));
 sky130_fd_sc_hd__a22o_2 _06231_ (.A1(\tag_array.tag0[9][4] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[10][4] ),
    .X(_03582_));
 sky130_fd_sc_hd__a221o_2 _06232_ (.A1(\tag_array.tag0[8][4] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[11][4] ),
    .C1(_03582_),
    .X(_03583_));
 sky130_fd_sc_hd__a22o_2 _06233_ (.A1(\tag_array.tag0[5][4] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[6][4] ),
    .X(_03584_));
 sky130_fd_sc_hd__a221o_2 _06234_ (.A1(\tag_array.tag0[4][4] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[7][4] ),
    .C1(_03584_),
    .X(_03585_));
 sky130_fd_sc_hd__a22o_2 _06235_ (.A1(\tag_array.tag0[13][4] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[14][4] ),
    .X(_03586_));
 sky130_fd_sc_hd__a221o_2 _06236_ (.A1(\tag_array.tag0[12][4] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[15][4] ),
    .C1(_03586_),
    .X(_03587_));
 sky130_fd_sc_hd__a22o_2 _06237_ (.A1(\tag_array.tag0[1][4] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[2][4] ),
    .X(_03588_));
 sky130_fd_sc_hd__a221o_2 _06238_ (.A1(\tag_array.tag0[0][4] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[3][4] ),
    .C1(_03588_),
    .X(_03589_));
 sky130_fd_sc_hd__a22o_2 _06239_ (.A1(_03506_),
    .A2(_03583_),
    .B1(_03587_),
    .B2(_03522_),
    .X(_03590_));
 sky130_fd_sc_hd__a22o_2 _06240_ (.A1(_03526_),
    .A2(_03585_),
    .B1(_03589_),
    .B2(_03518_),
    .X(_03591_));
 sky130_fd_sc_hd__or2_2 _06241_ (.A(_03590_),
    .B(_03591_),
    .X(_00150_));
 sky130_fd_sc_hd__a22o_2 _06242_ (.A1(\tag_array.tag0[13][5] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[14][5] ),
    .X(_03592_));
 sky130_fd_sc_hd__a221o_2 _06243_ (.A1(\tag_array.tag0[12][5] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[15][5] ),
    .C1(_03592_),
    .X(_03593_));
 sky130_fd_sc_hd__a22o_2 _06244_ (.A1(\tag_array.tag0[5][5] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[6][5] ),
    .X(_03594_));
 sky130_fd_sc_hd__a221o_2 _06245_ (.A1(\tag_array.tag0[4][5] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[7][5] ),
    .C1(_03594_),
    .X(_03595_));
 sky130_fd_sc_hd__a22o_2 _06246_ (.A1(\tag_array.tag0[9][5] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[10][5] ),
    .X(_03596_));
 sky130_fd_sc_hd__a221o_2 _06247_ (.A1(\tag_array.tag0[8][5] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[11][5] ),
    .C1(_03596_),
    .X(_03597_));
 sky130_fd_sc_hd__a22o_2 _06248_ (.A1(\tag_array.tag0[1][5] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[2][5] ),
    .X(_03598_));
 sky130_fd_sc_hd__a221o_2 _06249_ (.A1(\tag_array.tag0[0][5] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[3][5] ),
    .C1(_03598_),
    .X(_03599_));
 sky130_fd_sc_hd__a22o_2 _06250_ (.A1(_03522_),
    .A2(_03593_),
    .B1(_03597_),
    .B2(_03506_),
    .X(_03600_));
 sky130_fd_sc_hd__a22o_2 _06251_ (.A1(_03526_),
    .A2(_03595_),
    .B1(_03599_),
    .B2(_03518_),
    .X(_03601_));
 sky130_fd_sc_hd__or2_2 _06252_ (.A(_03600_),
    .B(_03601_),
    .X(_00151_));
 sky130_fd_sc_hd__a22o_2 _06253_ (.A1(\tag_array.tag0[13][6] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[14][6] ),
    .X(_03602_));
 sky130_fd_sc_hd__a221o_2 _06254_ (.A1(\tag_array.tag0[12][6] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[15][6] ),
    .C1(_03602_),
    .X(_03603_));
 sky130_fd_sc_hd__a22o_2 _06255_ (.A1(\tag_array.tag0[5][6] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[6][6] ),
    .X(_03604_));
 sky130_fd_sc_hd__a221o_2 _06256_ (.A1(\tag_array.tag0[4][6] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[7][6] ),
    .C1(_03604_),
    .X(_03605_));
 sky130_fd_sc_hd__a22o_2 _06257_ (.A1(\tag_array.tag0[9][6] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[10][6] ),
    .X(_03606_));
 sky130_fd_sc_hd__a221o_2 _06258_ (.A1(\tag_array.tag0[8][6] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[11][6] ),
    .C1(_03606_),
    .X(_03607_));
 sky130_fd_sc_hd__a22o_2 _06259_ (.A1(\tag_array.tag0[1][6] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[2][6] ),
    .X(_03608_));
 sky130_fd_sc_hd__a221o_2 _06260_ (.A1(\tag_array.tag0[0][6] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[3][6] ),
    .C1(_03608_),
    .X(_03609_));
 sky130_fd_sc_hd__a22o_2 _06261_ (.A1(_03522_),
    .A2(_03603_),
    .B1(_03607_),
    .B2(_03506_),
    .X(_03610_));
 sky130_fd_sc_hd__a22o_2 _06262_ (.A1(_03526_),
    .A2(_03605_),
    .B1(_03609_),
    .B2(_03518_),
    .X(_03611_));
 sky130_fd_sc_hd__or2_2 _06263_ (.A(_03610_),
    .B(_03611_),
    .X(_00152_));
 sky130_fd_sc_hd__a22o_2 _06264_ (.A1(\tag_array.tag0[9][7] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[10][7] ),
    .X(_03612_));
 sky130_fd_sc_hd__a221o_2 _06265_ (.A1(\tag_array.tag0[8][7] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[11][7] ),
    .C1(_03612_),
    .X(_03613_));
 sky130_fd_sc_hd__a22o_2 _06266_ (.A1(\tag_array.tag0[1][7] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[2][7] ),
    .X(_03614_));
 sky130_fd_sc_hd__a221o_2 _06267_ (.A1(\tag_array.tag0[0][7] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[3][7] ),
    .C1(_03614_),
    .X(_03615_));
 sky130_fd_sc_hd__a22o_2 _06268_ (.A1(\tag_array.tag0[13][7] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[14][7] ),
    .X(_03616_));
 sky130_fd_sc_hd__a221o_2 _06269_ (.A1(\tag_array.tag0[12][7] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[15][7] ),
    .C1(_03616_),
    .X(_03617_));
 sky130_fd_sc_hd__a22o_2 _06270_ (.A1(\tag_array.tag0[5][7] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[6][7] ),
    .X(_03618_));
 sky130_fd_sc_hd__a221o_2 _06271_ (.A1(\tag_array.tag0[4][7] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[7][7] ),
    .C1(_03618_),
    .X(_03619_));
 sky130_fd_sc_hd__a22o_2 _06272_ (.A1(_03506_),
    .A2(_03613_),
    .B1(_03617_),
    .B2(_03522_),
    .X(_03620_));
 sky130_fd_sc_hd__a22o_2 _06273_ (.A1(_03518_),
    .A2(_03615_),
    .B1(_03619_),
    .B2(_03526_),
    .X(_03621_));
 sky130_fd_sc_hd__or2_2 _06274_ (.A(_03620_),
    .B(_03621_),
    .X(_00153_));
 sky130_fd_sc_hd__a22o_2 _06275_ (.A1(\tag_array.tag0[9][8] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[10][8] ),
    .X(_03622_));
 sky130_fd_sc_hd__a221o_2 _06276_ (.A1(\tag_array.tag0[8][8] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[11][8] ),
    .C1(_03622_),
    .X(_03623_));
 sky130_fd_sc_hd__a22o_2 _06277_ (.A1(\tag_array.tag0[1][8] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[2][8] ),
    .X(_03624_));
 sky130_fd_sc_hd__a221o_2 _06278_ (.A1(\tag_array.tag0[0][8] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[3][8] ),
    .C1(_03624_),
    .X(_03625_));
 sky130_fd_sc_hd__a22o_2 _06279_ (.A1(\tag_array.tag0[13][8] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[14][8] ),
    .X(_03626_));
 sky130_fd_sc_hd__a221o_2 _06280_ (.A1(\tag_array.tag0[12][8] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[15][8] ),
    .C1(_03626_),
    .X(_03627_));
 sky130_fd_sc_hd__a22o_2 _06281_ (.A1(\tag_array.tag0[5][8] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[6][8] ),
    .X(_03628_));
 sky130_fd_sc_hd__a221o_2 _06282_ (.A1(\tag_array.tag0[4][8] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[7][8] ),
    .C1(_03628_),
    .X(_03629_));
 sky130_fd_sc_hd__a22o_2 _06283_ (.A1(_03506_),
    .A2(_03623_),
    .B1(_03627_),
    .B2(_03522_),
    .X(_03630_));
 sky130_fd_sc_hd__a22o_2 _06284_ (.A1(_03518_),
    .A2(_03625_),
    .B1(_03629_),
    .B2(_03526_),
    .X(_03631_));
 sky130_fd_sc_hd__or2_2 _06285_ (.A(_03630_),
    .B(_03631_),
    .X(_00154_));
 sky130_fd_sc_hd__a22o_2 _06286_ (.A1(\tag_array.tag0[13][9] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[14][9] ),
    .X(_03632_));
 sky130_fd_sc_hd__a221o_2 _06287_ (.A1(\tag_array.tag0[12][9] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[15][9] ),
    .C1(_03632_),
    .X(_03633_));
 sky130_fd_sc_hd__a22o_2 _06288_ (.A1(\tag_array.tag0[1][9] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[2][9] ),
    .X(_03634_));
 sky130_fd_sc_hd__a221o_2 _06289_ (.A1(\tag_array.tag0[0][9] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[3][9] ),
    .C1(_03634_),
    .X(_03635_));
 sky130_fd_sc_hd__a22o_2 _06290_ (.A1(\tag_array.tag0[9][9] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[10][9] ),
    .X(_03636_));
 sky130_fd_sc_hd__a221o_2 _06291_ (.A1(\tag_array.tag0[8][9] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[11][9] ),
    .C1(_03636_),
    .X(_03637_));
 sky130_fd_sc_hd__a22o_2 _06292_ (.A1(\tag_array.tag0[5][9] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[6][9] ),
    .X(_03638_));
 sky130_fd_sc_hd__a221o_2 _06293_ (.A1(\tag_array.tag0[4][9] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[7][9] ),
    .C1(_03638_),
    .X(_03639_));
 sky130_fd_sc_hd__a22o_2 _06294_ (.A1(_03522_),
    .A2(_03633_),
    .B1(_03637_),
    .B2(_03506_),
    .X(_03640_));
 sky130_fd_sc_hd__a22o_2 _06295_ (.A1(_03518_),
    .A2(_03635_),
    .B1(_03639_),
    .B2(_03526_),
    .X(_03641_));
 sky130_fd_sc_hd__or2_2 _06296_ (.A(_03640_),
    .B(_03641_),
    .X(_00155_));
 sky130_fd_sc_hd__a22o_2 _06297_ (.A1(\tag_array.tag0[13][10] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[14][10] ),
    .X(_03642_));
 sky130_fd_sc_hd__a221o_2 _06298_ (.A1(\tag_array.tag0[12][10] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[15][10] ),
    .C1(_03642_),
    .X(_03643_));
 sky130_fd_sc_hd__a22o_2 _06299_ (.A1(\tag_array.tag0[5][10] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[6][10] ),
    .X(_03644_));
 sky130_fd_sc_hd__a221o_2 _06300_ (.A1(\tag_array.tag0[4][10] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[7][10] ),
    .C1(_03644_),
    .X(_03645_));
 sky130_fd_sc_hd__a22o_2 _06301_ (.A1(\tag_array.tag0[9][10] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[10][10] ),
    .X(_03646_));
 sky130_fd_sc_hd__a221o_2 _06302_ (.A1(\tag_array.tag0[8][10] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[11][10] ),
    .C1(_03646_),
    .X(_03647_));
 sky130_fd_sc_hd__a22o_2 _06303_ (.A1(\tag_array.tag0[1][10] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[2][10] ),
    .X(_03648_));
 sky130_fd_sc_hd__a221o_2 _06304_ (.A1(\tag_array.tag0[0][10] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[3][10] ),
    .C1(_03648_),
    .X(_03649_));
 sky130_fd_sc_hd__a22o_2 _06305_ (.A1(_03522_),
    .A2(_03643_),
    .B1(_03647_),
    .B2(_03506_),
    .X(_03650_));
 sky130_fd_sc_hd__a22o_2 _06306_ (.A1(_03526_),
    .A2(_03645_),
    .B1(_03649_),
    .B2(_03518_),
    .X(_03651_));
 sky130_fd_sc_hd__or2_2 _06307_ (.A(_03650_),
    .B(_03651_),
    .X(_00132_));
 sky130_fd_sc_hd__a22o_2 _06308_ (.A1(\tag_array.tag0[13][11] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[14][11] ),
    .X(_03652_));
 sky130_fd_sc_hd__a221o_2 _06309_ (.A1(\tag_array.tag0[12][11] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[15][11] ),
    .C1(_03652_),
    .X(_03653_));
 sky130_fd_sc_hd__a22o_2 _06310_ (.A1(\tag_array.tag0[1][11] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[2][11] ),
    .X(_03654_));
 sky130_fd_sc_hd__a221o_2 _06311_ (.A1(\tag_array.tag0[0][11] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[3][11] ),
    .C1(_03654_),
    .X(_03655_));
 sky130_fd_sc_hd__a22o_2 _06312_ (.A1(\tag_array.tag0[9][11] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[10][11] ),
    .X(_03656_));
 sky130_fd_sc_hd__a221o_2 _06313_ (.A1(\tag_array.tag0[8][11] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[11][11] ),
    .C1(_03656_),
    .X(_03657_));
 sky130_fd_sc_hd__a22o_2 _06314_ (.A1(\tag_array.tag0[5][11] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[6][11] ),
    .X(_03658_));
 sky130_fd_sc_hd__a221o_2 _06315_ (.A1(\tag_array.tag0[4][11] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[7][11] ),
    .C1(_03658_),
    .X(_03659_));
 sky130_fd_sc_hd__a22o_2 _06316_ (.A1(_03522_),
    .A2(_03653_),
    .B1(_03657_),
    .B2(_03506_),
    .X(_03660_));
 sky130_fd_sc_hd__a22o_2 _06317_ (.A1(_03518_),
    .A2(_03655_),
    .B1(_03659_),
    .B2(_03526_),
    .X(_03661_));
 sky130_fd_sc_hd__or2_2 _06318_ (.A(_03660_),
    .B(_03661_),
    .X(_00133_));
 sky130_fd_sc_hd__a22o_2 _06319_ (.A1(\tag_array.tag0[9][12] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[10][12] ),
    .X(_03662_));
 sky130_fd_sc_hd__a221o_2 _06320_ (.A1(\tag_array.tag0[8][12] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[11][12] ),
    .C1(_03662_),
    .X(_03663_));
 sky130_fd_sc_hd__a22o_2 _06321_ (.A1(\tag_array.tag0[5][12] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[6][12] ),
    .X(_03664_));
 sky130_fd_sc_hd__a221o_2 _06322_ (.A1(\tag_array.tag0[4][12] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[7][12] ),
    .C1(_03664_),
    .X(_03665_));
 sky130_fd_sc_hd__a22o_2 _06323_ (.A1(\tag_array.tag0[13][12] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[14][12] ),
    .X(_03666_));
 sky130_fd_sc_hd__a221o_2 _06324_ (.A1(\tag_array.tag0[12][12] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[15][12] ),
    .C1(_03666_),
    .X(_03667_));
 sky130_fd_sc_hd__a22o_2 _06325_ (.A1(\tag_array.tag0[1][12] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[2][12] ),
    .X(_03668_));
 sky130_fd_sc_hd__a221o_2 _06326_ (.A1(\tag_array.tag0[0][12] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[3][12] ),
    .C1(_03668_),
    .X(_03669_));
 sky130_fd_sc_hd__a22o_2 _06327_ (.A1(_03506_),
    .A2(_03663_),
    .B1(_03667_),
    .B2(_03522_),
    .X(_03670_));
 sky130_fd_sc_hd__a22o_2 _06328_ (.A1(_03526_),
    .A2(_03665_),
    .B1(_03669_),
    .B2(_03518_),
    .X(_03671_));
 sky130_fd_sc_hd__or2_2 _06329_ (.A(_03670_),
    .B(_03671_),
    .X(_00134_));
 sky130_fd_sc_hd__a22o_2 _06330_ (.A1(\tag_array.tag0[9][13] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[10][13] ),
    .X(_03672_));
 sky130_fd_sc_hd__a221o_2 _06331_ (.A1(\tag_array.tag0[8][13] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[11][13] ),
    .C1(_03672_),
    .X(_03673_));
 sky130_fd_sc_hd__a22o_2 _06332_ (.A1(\tag_array.tag0[1][13] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[2][13] ),
    .X(_03674_));
 sky130_fd_sc_hd__a221o_2 _06333_ (.A1(\tag_array.tag0[0][13] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[3][13] ),
    .C1(_03674_),
    .X(_03675_));
 sky130_fd_sc_hd__a22o_2 _06334_ (.A1(\tag_array.tag0[13][13] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[14][13] ),
    .X(_03676_));
 sky130_fd_sc_hd__a221o_2 _06335_ (.A1(\tag_array.tag0[12][13] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[15][13] ),
    .C1(_03676_),
    .X(_03677_));
 sky130_fd_sc_hd__a22o_2 _06336_ (.A1(\tag_array.tag0[5][13] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[6][13] ),
    .X(_03678_));
 sky130_fd_sc_hd__a221o_2 _06337_ (.A1(\tag_array.tag0[4][13] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[7][13] ),
    .C1(_03678_),
    .X(_03679_));
 sky130_fd_sc_hd__a22o_2 _06338_ (.A1(_03506_),
    .A2(_03673_),
    .B1(_03677_),
    .B2(_03522_),
    .X(_03680_));
 sky130_fd_sc_hd__a22o_2 _06339_ (.A1(_03518_),
    .A2(_03675_),
    .B1(_03679_),
    .B2(_03526_),
    .X(_03681_));
 sky130_fd_sc_hd__or2_2 _06340_ (.A(_03680_),
    .B(_03681_),
    .X(_00135_));
 sky130_fd_sc_hd__a22o_2 _06341_ (.A1(\tag_array.tag0[9][14] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[10][14] ),
    .X(_03682_));
 sky130_fd_sc_hd__a221o_2 _06342_ (.A1(\tag_array.tag0[8][14] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[11][14] ),
    .C1(_03682_),
    .X(_03683_));
 sky130_fd_sc_hd__a22o_2 _06343_ (.A1(\tag_array.tag0[5][14] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[6][14] ),
    .X(_03684_));
 sky130_fd_sc_hd__a221o_2 _06344_ (.A1(\tag_array.tag0[4][14] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[7][14] ),
    .C1(_03684_),
    .X(_03685_));
 sky130_fd_sc_hd__a22o_2 _06345_ (.A1(\tag_array.tag0[13][14] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[14][14] ),
    .X(_03686_));
 sky130_fd_sc_hd__a221o_2 _06346_ (.A1(\tag_array.tag0[12][14] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[15][14] ),
    .C1(_03686_),
    .X(_03687_));
 sky130_fd_sc_hd__a22o_2 _06347_ (.A1(\tag_array.tag0[1][14] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[2][14] ),
    .X(_03688_));
 sky130_fd_sc_hd__a221o_2 _06348_ (.A1(\tag_array.tag0[0][14] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[3][14] ),
    .C1(_03688_),
    .X(_03689_));
 sky130_fd_sc_hd__a22o_2 _06349_ (.A1(_03506_),
    .A2(_03683_),
    .B1(_03687_),
    .B2(_03522_),
    .X(_03690_));
 sky130_fd_sc_hd__a22o_2 _06350_ (.A1(_03526_),
    .A2(_03685_),
    .B1(_03689_),
    .B2(_03518_),
    .X(_03691_));
 sky130_fd_sc_hd__or2_2 _06351_ (.A(_03690_),
    .B(_03691_),
    .X(_00136_));
 sky130_fd_sc_hd__a22o_2 _06352_ (.A1(\tag_array.tag0[13][15] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[14][15] ),
    .X(_03692_));
 sky130_fd_sc_hd__a221o_2 _06353_ (.A1(\tag_array.tag0[12][15] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[15][15] ),
    .C1(_03692_),
    .X(_03693_));
 sky130_fd_sc_hd__a22o_2 _06354_ (.A1(\tag_array.tag0[1][15] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[2][15] ),
    .X(_03694_));
 sky130_fd_sc_hd__a221o_2 _06355_ (.A1(\tag_array.tag0[0][15] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[3][15] ),
    .C1(_03694_),
    .X(_03695_));
 sky130_fd_sc_hd__a22o_2 _06356_ (.A1(\tag_array.tag0[9][15] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[10][15] ),
    .X(_03696_));
 sky130_fd_sc_hd__a221o_2 _06357_ (.A1(\tag_array.tag0[8][15] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[11][15] ),
    .C1(_03696_),
    .X(_03697_));
 sky130_fd_sc_hd__a22o_2 _06358_ (.A1(\tag_array.tag0[5][15] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[6][15] ),
    .X(_03698_));
 sky130_fd_sc_hd__a221o_2 _06359_ (.A1(\tag_array.tag0[4][15] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[7][15] ),
    .C1(_03698_),
    .X(_03699_));
 sky130_fd_sc_hd__a22o_2 _06360_ (.A1(_03522_),
    .A2(_03693_),
    .B1(_03697_),
    .B2(_03506_),
    .X(_03700_));
 sky130_fd_sc_hd__a22o_2 _06361_ (.A1(_03518_),
    .A2(_03695_),
    .B1(_03699_),
    .B2(_03526_),
    .X(_03701_));
 sky130_fd_sc_hd__or2_2 _06362_ (.A(_03700_),
    .B(_03701_),
    .X(_00137_));
 sky130_fd_sc_hd__a22o_2 _06363_ (.A1(\tag_array.tag0[9][16] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[10][16] ),
    .X(_03702_));
 sky130_fd_sc_hd__a221o_2 _06364_ (.A1(\tag_array.tag0[8][16] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[11][16] ),
    .C1(_03702_),
    .X(_03703_));
 sky130_fd_sc_hd__a22o_2 _06365_ (.A1(\tag_array.tag0[5][16] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[6][16] ),
    .X(_03704_));
 sky130_fd_sc_hd__a221o_2 _06366_ (.A1(\tag_array.tag0[4][16] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[7][16] ),
    .C1(_03704_),
    .X(_03705_));
 sky130_fd_sc_hd__a22o_2 _06367_ (.A1(\tag_array.tag0[13][16] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[14][16] ),
    .X(_03706_));
 sky130_fd_sc_hd__a221o_2 _06368_ (.A1(\tag_array.tag0[12][16] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[15][16] ),
    .C1(_03706_),
    .X(_03707_));
 sky130_fd_sc_hd__a22o_2 _06369_ (.A1(\tag_array.tag0[1][16] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[2][16] ),
    .X(_03708_));
 sky130_fd_sc_hd__a221o_2 _06370_ (.A1(\tag_array.tag0[0][16] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[3][16] ),
    .C1(_03708_),
    .X(_03709_));
 sky130_fd_sc_hd__a22o_2 _06371_ (.A1(_03506_),
    .A2(_03703_),
    .B1(_03707_),
    .B2(_03522_),
    .X(_03710_));
 sky130_fd_sc_hd__a22o_2 _06372_ (.A1(_03526_),
    .A2(_03705_),
    .B1(_03709_),
    .B2(_03518_),
    .X(_03711_));
 sky130_fd_sc_hd__or2_2 _06373_ (.A(_03710_),
    .B(_03711_),
    .X(_00138_));
 sky130_fd_sc_hd__a22o_2 _06374_ (.A1(\tag_array.tag0[13][17] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[14][17] ),
    .X(_03712_));
 sky130_fd_sc_hd__a221o_2 _06375_ (.A1(\tag_array.tag0[12][17] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[15][17] ),
    .C1(_03712_),
    .X(_03713_));
 sky130_fd_sc_hd__a22o_2 _06376_ (.A1(\tag_array.tag0[5][17] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[6][17] ),
    .X(_03714_));
 sky130_fd_sc_hd__a221o_2 _06377_ (.A1(\tag_array.tag0[4][17] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[7][17] ),
    .C1(_03714_),
    .X(_03715_));
 sky130_fd_sc_hd__a22o_2 _06378_ (.A1(\tag_array.tag0[9][17] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[10][17] ),
    .X(_03716_));
 sky130_fd_sc_hd__a221o_2 _06379_ (.A1(\tag_array.tag0[8][17] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[11][17] ),
    .C1(_03716_),
    .X(_03717_));
 sky130_fd_sc_hd__a22o_2 _06380_ (.A1(\tag_array.tag0[1][17] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[2][17] ),
    .X(_03718_));
 sky130_fd_sc_hd__a221o_2 _06381_ (.A1(\tag_array.tag0[0][17] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[3][17] ),
    .C1(_03718_),
    .X(_03719_));
 sky130_fd_sc_hd__a22o_2 _06382_ (.A1(_03522_),
    .A2(_03713_),
    .B1(_03717_),
    .B2(_03506_),
    .X(_03720_));
 sky130_fd_sc_hd__a22o_2 _06383_ (.A1(_03526_),
    .A2(_03715_),
    .B1(_03719_),
    .B2(_03518_),
    .X(_03721_));
 sky130_fd_sc_hd__or2_2 _06384_ (.A(_03720_),
    .B(_03721_),
    .X(_00139_));
 sky130_fd_sc_hd__a22o_2 _06385_ (.A1(\tag_array.tag0[13][18] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[14][18] ),
    .X(_03722_));
 sky130_fd_sc_hd__a221o_2 _06386_ (.A1(\tag_array.tag0[12][18] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[15][18] ),
    .C1(_03722_),
    .X(_03723_));
 sky130_fd_sc_hd__a22o_2 _06387_ (.A1(\tag_array.tag0[1][18] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[2][18] ),
    .X(_03724_));
 sky130_fd_sc_hd__a221o_2 _06388_ (.A1(\tag_array.tag0[0][18] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[3][18] ),
    .C1(_03724_),
    .X(_03725_));
 sky130_fd_sc_hd__a22o_2 _06389_ (.A1(\tag_array.tag0[9][18] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[10][18] ),
    .X(_03726_));
 sky130_fd_sc_hd__a221o_2 _06390_ (.A1(\tag_array.tag0[8][18] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[11][18] ),
    .C1(_03726_),
    .X(_03727_));
 sky130_fd_sc_hd__a22o_2 _06391_ (.A1(\tag_array.tag0[5][18] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[6][18] ),
    .X(_03728_));
 sky130_fd_sc_hd__a221o_2 _06392_ (.A1(\tag_array.tag0[4][18] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[7][18] ),
    .C1(_03728_),
    .X(_03729_));
 sky130_fd_sc_hd__a22o_2 _06393_ (.A1(_03522_),
    .A2(_03723_),
    .B1(_03727_),
    .B2(_03506_),
    .X(_03730_));
 sky130_fd_sc_hd__a22o_2 _06394_ (.A1(_03518_),
    .A2(_03725_),
    .B1(_03729_),
    .B2(_03526_),
    .X(_03731_));
 sky130_fd_sc_hd__or2_2 _06395_ (.A(_03730_),
    .B(_03731_),
    .X(_00140_));
 sky130_fd_sc_hd__a22o_2 _06396_ (.A1(\tag_array.tag0[13][19] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[14][19] ),
    .X(_03732_));
 sky130_fd_sc_hd__a221o_2 _06397_ (.A1(\tag_array.tag0[12][19] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[15][19] ),
    .C1(_03732_),
    .X(_03733_));
 sky130_fd_sc_hd__a22o_2 _06398_ (.A1(\tag_array.tag0[1][19] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[2][19] ),
    .X(_03734_));
 sky130_fd_sc_hd__a221o_2 _06399_ (.A1(\tag_array.tag0[0][19] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[3][19] ),
    .C1(_03734_),
    .X(_03735_));
 sky130_fd_sc_hd__a22o_2 _06400_ (.A1(\tag_array.tag0[9][19] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[10][19] ),
    .X(_03736_));
 sky130_fd_sc_hd__a221o_2 _06401_ (.A1(\tag_array.tag0[8][19] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[11][19] ),
    .C1(_03736_),
    .X(_03737_));
 sky130_fd_sc_hd__a22o_2 _06402_ (.A1(\tag_array.tag0[5][19] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[6][19] ),
    .X(_03738_));
 sky130_fd_sc_hd__a221o_2 _06403_ (.A1(\tag_array.tag0[4][19] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[7][19] ),
    .C1(_03738_),
    .X(_03739_));
 sky130_fd_sc_hd__a22o_2 _06404_ (.A1(_03522_),
    .A2(_03733_),
    .B1(_03737_),
    .B2(_03506_),
    .X(_03740_));
 sky130_fd_sc_hd__a22o_2 _06405_ (.A1(_03518_),
    .A2(_03735_),
    .B1(_03739_),
    .B2(_03526_),
    .X(_03741_));
 sky130_fd_sc_hd__or2_2 _06406_ (.A(_03740_),
    .B(_03741_),
    .X(_00141_));
 sky130_fd_sc_hd__a22o_2 _06407_ (.A1(\tag_array.tag0[13][20] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[14][20] ),
    .X(_03742_));
 sky130_fd_sc_hd__a221o_2 _06408_ (.A1(\tag_array.tag0[12][20] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[15][20] ),
    .C1(_03742_),
    .X(_03743_));
 sky130_fd_sc_hd__a22o_2 _06409_ (.A1(\tag_array.tag0[5][20] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[6][20] ),
    .X(_03744_));
 sky130_fd_sc_hd__a221o_2 _06410_ (.A1(\tag_array.tag0[4][20] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[7][20] ),
    .C1(_03744_),
    .X(_03745_));
 sky130_fd_sc_hd__a22o_2 _06411_ (.A1(\tag_array.tag0[9][20] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[10][20] ),
    .X(_03746_));
 sky130_fd_sc_hd__a221o_2 _06412_ (.A1(\tag_array.tag0[8][20] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[11][20] ),
    .C1(_03746_),
    .X(_03747_));
 sky130_fd_sc_hd__a22o_2 _06413_ (.A1(\tag_array.tag0[1][20] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[2][20] ),
    .X(_03748_));
 sky130_fd_sc_hd__a221o_2 _06414_ (.A1(\tag_array.tag0[0][20] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[3][20] ),
    .C1(_03748_),
    .X(_03749_));
 sky130_fd_sc_hd__a22o_2 _06415_ (.A1(_03522_),
    .A2(_03743_),
    .B1(_03747_),
    .B2(_03506_),
    .X(_03750_));
 sky130_fd_sc_hd__a22o_2 _06416_ (.A1(_03526_),
    .A2(_03745_),
    .B1(_03749_),
    .B2(_03518_),
    .X(_03751_));
 sky130_fd_sc_hd__or2_2 _06417_ (.A(_03750_),
    .B(_03751_),
    .X(_00143_));
 sky130_fd_sc_hd__a22o_2 _06418_ (.A1(\tag_array.tag0[13][21] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[14][21] ),
    .X(_03752_));
 sky130_fd_sc_hd__a221o_2 _06419_ (.A1(\tag_array.tag0[12][21] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[15][21] ),
    .C1(_03752_),
    .X(_03753_));
 sky130_fd_sc_hd__a22o_2 _06420_ (.A1(\tag_array.tag0[5][21] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[6][21] ),
    .X(_03754_));
 sky130_fd_sc_hd__a221o_2 _06421_ (.A1(\tag_array.tag0[4][21] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[7][21] ),
    .C1(_03754_),
    .X(_03755_));
 sky130_fd_sc_hd__a22o_2 _06422_ (.A1(\tag_array.tag0[9][21] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[10][21] ),
    .X(_03756_));
 sky130_fd_sc_hd__a221o_2 _06423_ (.A1(\tag_array.tag0[8][21] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[11][21] ),
    .C1(_03756_),
    .X(_03757_));
 sky130_fd_sc_hd__a22o_2 _06424_ (.A1(\tag_array.tag0[1][21] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[2][21] ),
    .X(_03758_));
 sky130_fd_sc_hd__a221o_2 _06425_ (.A1(\tag_array.tag0[0][21] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[3][21] ),
    .C1(_03758_),
    .X(_03759_));
 sky130_fd_sc_hd__a22o_2 _06426_ (.A1(_03522_),
    .A2(_03753_),
    .B1(_03757_),
    .B2(_03506_),
    .X(_03760_));
 sky130_fd_sc_hd__a22o_2 _06427_ (.A1(_03526_),
    .A2(_03755_),
    .B1(_03759_),
    .B2(_03518_),
    .X(_03761_));
 sky130_fd_sc_hd__or2_2 _06428_ (.A(_03760_),
    .B(_03761_),
    .X(_00144_));
 sky130_fd_sc_hd__a22o_2 _06429_ (.A1(\tag_array.tag0[9][22] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[10][22] ),
    .X(_03762_));
 sky130_fd_sc_hd__a221o_2 _06430_ (.A1(\tag_array.tag0[8][22] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[11][22] ),
    .C1(_03762_),
    .X(_03763_));
 sky130_fd_sc_hd__a22o_2 _06431_ (.A1(\tag_array.tag0[5][22] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[6][22] ),
    .X(_03764_));
 sky130_fd_sc_hd__a221o_2 _06432_ (.A1(\tag_array.tag0[4][22] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[7][22] ),
    .C1(_03764_),
    .X(_03765_));
 sky130_fd_sc_hd__a22o_2 _06433_ (.A1(\tag_array.tag0[13][22] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[14][22] ),
    .X(_03766_));
 sky130_fd_sc_hd__a221o_2 _06434_ (.A1(\tag_array.tag0[12][22] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[15][22] ),
    .C1(_03766_),
    .X(_03767_));
 sky130_fd_sc_hd__a22o_2 _06435_ (.A1(\tag_array.tag0[1][22] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[2][22] ),
    .X(_03768_));
 sky130_fd_sc_hd__a221o_2 _06436_ (.A1(\tag_array.tag0[0][22] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[3][22] ),
    .C1(_03768_),
    .X(_03769_));
 sky130_fd_sc_hd__a22o_2 _06437_ (.A1(_03506_),
    .A2(_03763_),
    .B1(_03767_),
    .B2(_03522_),
    .X(_03770_));
 sky130_fd_sc_hd__a22o_2 _06438_ (.A1(_03526_),
    .A2(_03765_),
    .B1(_03769_),
    .B2(_03518_),
    .X(_03771_));
 sky130_fd_sc_hd__or2_2 _06439_ (.A(_03770_),
    .B(_03771_),
    .X(_00145_));
 sky130_fd_sc_hd__a22o_2 _06440_ (.A1(\tag_array.tag0[9][23] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[10][23] ),
    .X(_03772_));
 sky130_fd_sc_hd__a221o_2 _06441_ (.A1(\tag_array.tag0[8][23] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[11][23] ),
    .C1(_03772_),
    .X(_03773_));
 sky130_fd_sc_hd__a22o_2 _06442_ (.A1(\tag_array.tag0[1][23] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[2][23] ),
    .X(_03774_));
 sky130_fd_sc_hd__a221o_2 _06443_ (.A1(\tag_array.tag0[0][23] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[3][23] ),
    .C1(_03774_),
    .X(_03775_));
 sky130_fd_sc_hd__a22o_2 _06444_ (.A1(\tag_array.tag0[13][23] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[14][23] ),
    .X(_03776_));
 sky130_fd_sc_hd__a221o_2 _06445_ (.A1(\tag_array.tag0[12][23] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[15][23] ),
    .C1(_03776_),
    .X(_03777_));
 sky130_fd_sc_hd__a22o_2 _06446_ (.A1(\tag_array.tag0[5][23] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[6][23] ),
    .X(_03778_));
 sky130_fd_sc_hd__a221o_2 _06447_ (.A1(\tag_array.tag0[4][23] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[7][23] ),
    .C1(_03778_),
    .X(_03779_));
 sky130_fd_sc_hd__a22o_2 _06448_ (.A1(_03506_),
    .A2(_03773_),
    .B1(_03777_),
    .B2(_03522_),
    .X(_03780_));
 sky130_fd_sc_hd__a22o_2 _06449_ (.A1(_03518_),
    .A2(_03775_),
    .B1(_03779_),
    .B2(_03526_),
    .X(_03781_));
 sky130_fd_sc_hd__or2_2 _06450_ (.A(_03780_),
    .B(_03781_),
    .X(_00146_));
 sky130_fd_sc_hd__a22o_2 _06451_ (.A1(\tag_array.tag0[9][24] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[10][24] ),
    .X(_03782_));
 sky130_fd_sc_hd__a221o_2 _06452_ (.A1(\tag_array.tag0[8][24] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[11][24] ),
    .C1(_03782_),
    .X(_03783_));
 sky130_fd_sc_hd__a22o_2 _06453_ (.A1(\tag_array.tag0[1][24] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[2][24] ),
    .X(_03784_));
 sky130_fd_sc_hd__a221o_2 _06454_ (.A1(\tag_array.tag0[0][24] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[3][24] ),
    .C1(_03784_),
    .X(_03785_));
 sky130_fd_sc_hd__a22o_2 _06455_ (.A1(\tag_array.tag0[13][24] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[14][24] ),
    .X(_03786_));
 sky130_fd_sc_hd__a221o_2 _06456_ (.A1(\tag_array.tag0[12][24] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[15][24] ),
    .C1(_03786_),
    .X(_03787_));
 sky130_fd_sc_hd__a22o_2 _06457_ (.A1(\tag_array.tag0[5][24] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag0[6][24] ),
    .X(_03788_));
 sky130_fd_sc_hd__a221o_2 _06458_ (.A1(\tag_array.tag0[4][24] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag0[7][24] ),
    .C1(_03788_),
    .X(_03789_));
 sky130_fd_sc_hd__a22o_2 _06459_ (.A1(_03506_),
    .A2(_03783_),
    .B1(_03787_),
    .B2(_03522_),
    .X(_03790_));
 sky130_fd_sc_hd__a22o_2 _06460_ (.A1(_03518_),
    .A2(_03785_),
    .B1(_03789_),
    .B2(_03526_),
    .X(_03791_));
 sky130_fd_sc_hd__or2_2 _06461_ (.A(_03790_),
    .B(_03791_),
    .X(_00147_));
 sky130_fd_sc_hd__a22o_2 _06462_ (.A1(\tag_array.tag1[9][0] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[10][0] ),
    .X(_03792_));
 sky130_fd_sc_hd__a221o_2 _06463_ (.A1(\tag_array.tag1[8][0] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[11][0] ),
    .C1(_03792_),
    .X(_03793_));
 sky130_fd_sc_hd__a22o_2 _06464_ (.A1(\tag_array.tag1[1][0] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[2][0] ),
    .X(_03794_));
 sky130_fd_sc_hd__a221o_2 _06465_ (.A1(\tag_array.tag1[0][0] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[3][0] ),
    .C1(_03794_),
    .X(_03795_));
 sky130_fd_sc_hd__a22o_2 _06466_ (.A1(\tag_array.tag1[13][0] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[14][0] ),
    .X(_03796_));
 sky130_fd_sc_hd__a221o_2 _06467_ (.A1(\tag_array.tag1[12][0] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[15][0] ),
    .C1(_03796_),
    .X(_03797_));
 sky130_fd_sc_hd__a22o_2 _06468_ (.A1(\tag_array.tag1[5][0] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[6][0] ),
    .X(_03798_));
 sky130_fd_sc_hd__a221o_2 _06469_ (.A1(\tag_array.tag1[4][0] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[7][0] ),
    .C1(_03798_),
    .X(_03799_));
 sky130_fd_sc_hd__a22o_2 _06470_ (.A1(_03506_),
    .A2(_03793_),
    .B1(_03797_),
    .B2(_03522_),
    .X(_03800_));
 sky130_fd_sc_hd__a22o_2 _06471_ (.A1(_03518_),
    .A2(_03795_),
    .B1(_03799_),
    .B2(_03526_),
    .X(_03801_));
 sky130_fd_sc_hd__or2_2 _06472_ (.A(_03800_),
    .B(_03801_),
    .X(_00156_));
 sky130_fd_sc_hd__a22o_2 _06473_ (.A1(\tag_array.tag1[13][1] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[14][1] ),
    .X(_03802_));
 sky130_fd_sc_hd__a221o_2 _06474_ (.A1(\tag_array.tag1[12][1] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[15][1] ),
    .C1(_03802_),
    .X(_03803_));
 sky130_fd_sc_hd__a22o_2 _06475_ (.A1(\tag_array.tag1[5][1] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[6][1] ),
    .X(_03804_));
 sky130_fd_sc_hd__a221o_2 _06476_ (.A1(\tag_array.tag1[4][1] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[7][1] ),
    .C1(_03804_),
    .X(_03805_));
 sky130_fd_sc_hd__a22o_2 _06477_ (.A1(\tag_array.tag1[9][1] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[10][1] ),
    .X(_03806_));
 sky130_fd_sc_hd__a221o_2 _06478_ (.A1(\tag_array.tag1[8][1] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[11][1] ),
    .C1(_03806_),
    .X(_03807_));
 sky130_fd_sc_hd__a22o_2 _06479_ (.A1(\tag_array.tag1[1][1] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[2][1] ),
    .X(_03808_));
 sky130_fd_sc_hd__a221o_2 _06480_ (.A1(\tag_array.tag1[0][1] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[3][1] ),
    .C1(_03808_),
    .X(_03809_));
 sky130_fd_sc_hd__a22o_2 _06481_ (.A1(_03522_),
    .A2(_03803_),
    .B1(_03807_),
    .B2(_03506_),
    .X(_03810_));
 sky130_fd_sc_hd__a22o_2 _06482_ (.A1(_03526_),
    .A2(_03805_),
    .B1(_03809_),
    .B2(_03518_),
    .X(_03811_));
 sky130_fd_sc_hd__or2_2 _06483_ (.A(_03810_),
    .B(_03811_),
    .X(_00167_));
 sky130_fd_sc_hd__a22o_2 _06484_ (.A1(\tag_array.tag1[9][2] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[10][2] ),
    .X(_03812_));
 sky130_fd_sc_hd__a221o_2 _06485_ (.A1(\tag_array.tag1[8][2] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[11][2] ),
    .C1(_03812_),
    .X(_03813_));
 sky130_fd_sc_hd__a22o_2 _06486_ (.A1(\tag_array.tag1[5][2] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[6][2] ),
    .X(_03814_));
 sky130_fd_sc_hd__a221o_2 _06487_ (.A1(\tag_array.tag1[4][2] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[7][2] ),
    .C1(_03814_),
    .X(_03815_));
 sky130_fd_sc_hd__a22o_2 _06488_ (.A1(\tag_array.tag1[13][2] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[14][2] ),
    .X(_03816_));
 sky130_fd_sc_hd__a221o_2 _06489_ (.A1(\tag_array.tag1[12][2] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[15][2] ),
    .C1(_03816_),
    .X(_03817_));
 sky130_fd_sc_hd__a22o_2 _06490_ (.A1(\tag_array.tag1[1][2] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[2][2] ),
    .X(_03818_));
 sky130_fd_sc_hd__a221o_2 _06491_ (.A1(\tag_array.tag1[0][2] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[3][2] ),
    .C1(_03818_),
    .X(_03819_));
 sky130_fd_sc_hd__a22o_2 _06492_ (.A1(_03506_),
    .A2(_03813_),
    .B1(_03817_),
    .B2(_03522_),
    .X(_03820_));
 sky130_fd_sc_hd__a22o_2 _06493_ (.A1(_03526_),
    .A2(_03815_),
    .B1(_03819_),
    .B2(_03518_),
    .X(_03821_));
 sky130_fd_sc_hd__or2_2 _06494_ (.A(_03820_),
    .B(_03821_),
    .X(_00173_));
 sky130_fd_sc_hd__a22o_2 _06495_ (.A1(\tag_array.tag1[9][3] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[10][3] ),
    .X(_03822_));
 sky130_fd_sc_hd__a221o_2 _06496_ (.A1(\tag_array.tag1[8][3] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[11][3] ),
    .C1(_03822_),
    .X(_03823_));
 sky130_fd_sc_hd__a22o_2 _06497_ (.A1(\tag_array.tag1[5][3] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[6][3] ),
    .X(_03824_));
 sky130_fd_sc_hd__a221o_2 _06498_ (.A1(\tag_array.tag1[4][3] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[7][3] ),
    .C1(_03824_),
    .X(_03825_));
 sky130_fd_sc_hd__a22o_2 _06499_ (.A1(\tag_array.tag1[13][3] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[14][3] ),
    .X(_03826_));
 sky130_fd_sc_hd__a221o_2 _06500_ (.A1(\tag_array.tag1[12][3] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[15][3] ),
    .C1(_03826_),
    .X(_03827_));
 sky130_fd_sc_hd__a22o_2 _06501_ (.A1(\tag_array.tag1[1][3] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[2][3] ),
    .X(_03828_));
 sky130_fd_sc_hd__a221o_2 _06502_ (.A1(\tag_array.tag1[0][3] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[3][3] ),
    .C1(_03828_),
    .X(_03829_));
 sky130_fd_sc_hd__a22o_2 _06503_ (.A1(_03506_),
    .A2(_03823_),
    .B1(_03827_),
    .B2(_03522_),
    .X(_03830_));
 sky130_fd_sc_hd__a22o_2 _06504_ (.A1(_03526_),
    .A2(_03825_),
    .B1(_03829_),
    .B2(_03518_),
    .X(_03831_));
 sky130_fd_sc_hd__or2_2 _06505_ (.A(_03830_),
    .B(_03831_),
    .X(_00174_));
 sky130_fd_sc_hd__a22o_2 _06506_ (.A1(\tag_array.tag1[9][4] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[10][4] ),
    .X(_03832_));
 sky130_fd_sc_hd__a221o_2 _06507_ (.A1(\tag_array.tag1[8][4] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[11][4] ),
    .C1(_03832_),
    .X(_03833_));
 sky130_fd_sc_hd__a22o_2 _06508_ (.A1(\tag_array.tag1[1][4] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[2][4] ),
    .X(_03834_));
 sky130_fd_sc_hd__a221o_2 _06509_ (.A1(\tag_array.tag1[0][4] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[3][4] ),
    .C1(_03834_),
    .X(_03835_));
 sky130_fd_sc_hd__a22o_2 _06510_ (.A1(\tag_array.tag1[13][4] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[14][4] ),
    .X(_03836_));
 sky130_fd_sc_hd__a221o_2 _06511_ (.A1(\tag_array.tag1[12][4] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[15][4] ),
    .C1(_03836_),
    .X(_03837_));
 sky130_fd_sc_hd__a22o_2 _06512_ (.A1(\tag_array.tag1[5][4] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[6][4] ),
    .X(_03838_));
 sky130_fd_sc_hd__a221o_2 _06513_ (.A1(\tag_array.tag1[4][4] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[7][4] ),
    .C1(_03838_),
    .X(_03839_));
 sky130_fd_sc_hd__a22o_2 _06514_ (.A1(_03506_),
    .A2(_03833_),
    .B1(_03837_),
    .B2(_03522_),
    .X(_03840_));
 sky130_fd_sc_hd__a22o_2 _06515_ (.A1(_03518_),
    .A2(_03835_),
    .B1(_03839_),
    .B2(_03526_),
    .X(_03841_));
 sky130_fd_sc_hd__or2_2 _06516_ (.A(_03840_),
    .B(_03841_),
    .X(_00175_));
 sky130_fd_sc_hd__a22o_2 _06517_ (.A1(\tag_array.tag1[9][5] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[10][5] ),
    .X(_03842_));
 sky130_fd_sc_hd__a221o_2 _06518_ (.A1(\tag_array.tag1[8][5] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[11][5] ),
    .C1(_03842_),
    .X(_03843_));
 sky130_fd_sc_hd__a22o_2 _06519_ (.A1(\tag_array.tag1[1][5] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[2][5] ),
    .X(_03844_));
 sky130_fd_sc_hd__a221o_2 _06520_ (.A1(\tag_array.tag1[0][5] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[3][5] ),
    .C1(_03844_),
    .X(_03845_));
 sky130_fd_sc_hd__a22o_2 _06521_ (.A1(\tag_array.tag1[13][5] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[14][5] ),
    .X(_03846_));
 sky130_fd_sc_hd__a221o_2 _06522_ (.A1(\tag_array.tag1[12][5] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[15][5] ),
    .C1(_03846_),
    .X(_03847_));
 sky130_fd_sc_hd__a22o_2 _06523_ (.A1(\tag_array.tag1[5][5] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[6][5] ),
    .X(_03848_));
 sky130_fd_sc_hd__a221o_2 _06524_ (.A1(\tag_array.tag1[4][5] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[7][5] ),
    .C1(_03848_),
    .X(_03849_));
 sky130_fd_sc_hd__a22o_2 _06525_ (.A1(_03506_),
    .A2(_03843_),
    .B1(_03847_),
    .B2(_03522_),
    .X(_03850_));
 sky130_fd_sc_hd__a22o_2 _06526_ (.A1(_03518_),
    .A2(_03845_),
    .B1(_03849_),
    .B2(_03526_),
    .X(_03851_));
 sky130_fd_sc_hd__or2_2 _06527_ (.A(_03850_),
    .B(_03851_),
    .X(_00176_));
 sky130_fd_sc_hd__a22o_2 _06528_ (.A1(\tag_array.tag1[13][6] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[14][6] ),
    .X(_03852_));
 sky130_fd_sc_hd__a221o_2 _06529_ (.A1(\tag_array.tag1[12][6] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[15][6] ),
    .C1(_03852_),
    .X(_03853_));
 sky130_fd_sc_hd__a22o_2 _06530_ (.A1(\tag_array.tag1[1][6] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[2][6] ),
    .X(_03854_));
 sky130_fd_sc_hd__a221o_2 _06531_ (.A1(\tag_array.tag1[0][6] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[3][6] ),
    .C1(_03854_),
    .X(_03855_));
 sky130_fd_sc_hd__a22o_2 _06532_ (.A1(\tag_array.tag1[9][6] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[10][6] ),
    .X(_03856_));
 sky130_fd_sc_hd__a221o_2 _06533_ (.A1(\tag_array.tag1[8][6] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[11][6] ),
    .C1(_03856_),
    .X(_03857_));
 sky130_fd_sc_hd__a22o_2 _06534_ (.A1(\tag_array.tag1[5][6] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[6][6] ),
    .X(_03858_));
 sky130_fd_sc_hd__a221o_2 _06535_ (.A1(\tag_array.tag1[4][6] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[7][6] ),
    .C1(_03858_),
    .X(_03859_));
 sky130_fd_sc_hd__a22o_2 _06536_ (.A1(_03522_),
    .A2(_03853_),
    .B1(_03857_),
    .B2(_03506_),
    .X(_03860_));
 sky130_fd_sc_hd__a22o_2 _06537_ (.A1(_03518_),
    .A2(_03855_),
    .B1(_03859_),
    .B2(_03526_),
    .X(_03861_));
 sky130_fd_sc_hd__or2_2 _06538_ (.A(_03860_),
    .B(_03861_),
    .X(_00177_));
 sky130_fd_sc_hd__a22o_2 _06539_ (.A1(\tag_array.tag1[9][7] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[10][7] ),
    .X(_03862_));
 sky130_fd_sc_hd__a221o_2 _06540_ (.A1(\tag_array.tag1[8][7] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[11][7] ),
    .C1(_03862_),
    .X(_03863_));
 sky130_fd_sc_hd__a22o_2 _06541_ (.A1(\tag_array.tag1[5][7] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[6][7] ),
    .X(_03864_));
 sky130_fd_sc_hd__a221o_2 _06542_ (.A1(\tag_array.tag1[4][7] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[7][7] ),
    .C1(_03864_),
    .X(_03865_));
 sky130_fd_sc_hd__a22o_2 _06543_ (.A1(\tag_array.tag1[13][7] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[14][7] ),
    .X(_03866_));
 sky130_fd_sc_hd__a221o_2 _06544_ (.A1(\tag_array.tag1[12][7] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[15][7] ),
    .C1(_03866_),
    .X(_03867_));
 sky130_fd_sc_hd__a22o_2 _06545_ (.A1(\tag_array.tag1[1][7] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[2][7] ),
    .X(_03868_));
 sky130_fd_sc_hd__a221o_2 _06546_ (.A1(\tag_array.tag1[0][7] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[3][7] ),
    .C1(_03868_),
    .X(_03869_));
 sky130_fd_sc_hd__a22o_2 _06547_ (.A1(_03506_),
    .A2(_03863_),
    .B1(_03867_),
    .B2(_03522_),
    .X(_03870_));
 sky130_fd_sc_hd__a22o_2 _06548_ (.A1(_03526_),
    .A2(_03865_),
    .B1(_03869_),
    .B2(_03518_),
    .X(_03871_));
 sky130_fd_sc_hd__or2_2 _06549_ (.A(_03870_),
    .B(_03871_),
    .X(_00178_));
 sky130_fd_sc_hd__a22o_2 _06550_ (.A1(\tag_array.tag1[9][8] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[10][8] ),
    .X(_03872_));
 sky130_fd_sc_hd__a221o_2 _06551_ (.A1(\tag_array.tag1[8][8] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[11][8] ),
    .C1(_03872_),
    .X(_03873_));
 sky130_fd_sc_hd__a22o_2 _06552_ (.A1(\tag_array.tag1[5][8] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[6][8] ),
    .X(_03874_));
 sky130_fd_sc_hd__a221o_2 _06553_ (.A1(\tag_array.tag1[4][8] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[7][8] ),
    .C1(_03874_),
    .X(_03875_));
 sky130_fd_sc_hd__a22o_2 _06554_ (.A1(\tag_array.tag1[13][8] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[14][8] ),
    .X(_03876_));
 sky130_fd_sc_hd__a221o_2 _06555_ (.A1(\tag_array.tag1[12][8] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[15][8] ),
    .C1(_03876_),
    .X(_03877_));
 sky130_fd_sc_hd__a22o_2 _06556_ (.A1(\tag_array.tag1[1][8] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[2][8] ),
    .X(_03878_));
 sky130_fd_sc_hd__a221o_2 _06557_ (.A1(\tag_array.tag1[0][8] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[3][8] ),
    .C1(_03878_),
    .X(_03879_));
 sky130_fd_sc_hd__a22o_2 _06558_ (.A1(_03506_),
    .A2(_03873_),
    .B1(_03877_),
    .B2(_03522_),
    .X(_03880_));
 sky130_fd_sc_hd__a22o_2 _06559_ (.A1(_03526_),
    .A2(_03875_),
    .B1(_03879_),
    .B2(_03518_),
    .X(_03881_));
 sky130_fd_sc_hd__or2_2 _06560_ (.A(_03880_),
    .B(_03881_),
    .X(_00179_));
 sky130_fd_sc_hd__a22o_2 _06561_ (.A1(\tag_array.tag1[9][9] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[10][9] ),
    .X(_03882_));
 sky130_fd_sc_hd__a221o_2 _06562_ (.A1(\tag_array.tag1[8][9] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[11][9] ),
    .C1(_03882_),
    .X(_03883_));
 sky130_fd_sc_hd__a22o_2 _06563_ (.A1(\tag_array.tag1[5][9] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[6][9] ),
    .X(_03884_));
 sky130_fd_sc_hd__a221o_2 _06564_ (.A1(\tag_array.tag1[4][9] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[7][9] ),
    .C1(_03884_),
    .X(_03885_));
 sky130_fd_sc_hd__a22o_2 _06565_ (.A1(\tag_array.tag1[13][9] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[14][9] ),
    .X(_03886_));
 sky130_fd_sc_hd__a221o_2 _06566_ (.A1(\tag_array.tag1[12][9] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[15][9] ),
    .C1(_03886_),
    .X(_03887_));
 sky130_fd_sc_hd__a22o_2 _06567_ (.A1(\tag_array.tag1[1][9] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[2][9] ),
    .X(_03888_));
 sky130_fd_sc_hd__a221o_2 _06568_ (.A1(\tag_array.tag1[0][9] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[3][9] ),
    .C1(_03888_),
    .X(_03889_));
 sky130_fd_sc_hd__a22o_2 _06569_ (.A1(_03506_),
    .A2(_03883_),
    .B1(_03887_),
    .B2(_03522_),
    .X(_03890_));
 sky130_fd_sc_hd__a22o_2 _06570_ (.A1(_03526_),
    .A2(_03885_),
    .B1(_03889_),
    .B2(_03518_),
    .X(_03891_));
 sky130_fd_sc_hd__or2_2 _06571_ (.A(_03890_),
    .B(_03891_),
    .X(_00180_));
 sky130_fd_sc_hd__a22o_2 _06572_ (.A1(\tag_array.tag1[13][10] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[14][10] ),
    .X(_03892_));
 sky130_fd_sc_hd__a221o_2 _06573_ (.A1(\tag_array.tag1[12][10] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[15][10] ),
    .C1(_03892_),
    .X(_03893_));
 sky130_fd_sc_hd__a22o_2 _06574_ (.A1(\tag_array.tag1[1][10] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[2][10] ),
    .X(_03894_));
 sky130_fd_sc_hd__a221o_2 _06575_ (.A1(\tag_array.tag1[0][10] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[3][10] ),
    .C1(_03894_),
    .X(_03895_));
 sky130_fd_sc_hd__a22o_2 _06576_ (.A1(\tag_array.tag1[9][10] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[10][10] ),
    .X(_03896_));
 sky130_fd_sc_hd__a221o_2 _06577_ (.A1(\tag_array.tag1[8][10] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[11][10] ),
    .C1(_03896_),
    .X(_03897_));
 sky130_fd_sc_hd__a22o_2 _06578_ (.A1(\tag_array.tag1[5][10] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[6][10] ),
    .X(_03898_));
 sky130_fd_sc_hd__a221o_2 _06579_ (.A1(\tag_array.tag1[4][10] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[7][10] ),
    .C1(_03898_),
    .X(_03899_));
 sky130_fd_sc_hd__a22o_2 _06580_ (.A1(_03522_),
    .A2(_03893_),
    .B1(_03897_),
    .B2(_03506_),
    .X(_03900_));
 sky130_fd_sc_hd__a22o_2 _06581_ (.A1(_03518_),
    .A2(_03895_),
    .B1(_03899_),
    .B2(_03526_),
    .X(_03901_));
 sky130_fd_sc_hd__or2_2 _06582_ (.A(_03900_),
    .B(_03901_),
    .X(_00157_));
 sky130_fd_sc_hd__a22o_2 _06583_ (.A1(\tag_array.tag1[9][11] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[10][11] ),
    .X(_03902_));
 sky130_fd_sc_hd__a221o_2 _06584_ (.A1(\tag_array.tag1[8][11] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[11][11] ),
    .C1(_03902_),
    .X(_03903_));
 sky130_fd_sc_hd__a22o_2 _06585_ (.A1(\tag_array.tag1[5][11] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[6][11] ),
    .X(_03904_));
 sky130_fd_sc_hd__a221o_2 _06586_ (.A1(\tag_array.tag1[4][11] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[7][11] ),
    .C1(_03904_),
    .X(_03905_));
 sky130_fd_sc_hd__a22o_2 _06587_ (.A1(\tag_array.tag1[13][11] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[14][11] ),
    .X(_03906_));
 sky130_fd_sc_hd__a221o_2 _06588_ (.A1(\tag_array.tag1[12][11] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[15][11] ),
    .C1(_03906_),
    .X(_03907_));
 sky130_fd_sc_hd__a22o_2 _06589_ (.A1(\tag_array.tag1[1][11] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[2][11] ),
    .X(_03908_));
 sky130_fd_sc_hd__a221o_2 _06590_ (.A1(\tag_array.tag1[0][11] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[3][11] ),
    .C1(_03908_),
    .X(_03909_));
 sky130_fd_sc_hd__a22o_2 _06591_ (.A1(_03506_),
    .A2(_03903_),
    .B1(_03907_),
    .B2(_03522_),
    .X(_03910_));
 sky130_fd_sc_hd__a22o_2 _06592_ (.A1(_03526_),
    .A2(_03905_),
    .B1(_03909_),
    .B2(_03518_),
    .X(_03911_));
 sky130_fd_sc_hd__or2_2 _06593_ (.A(_03910_),
    .B(_03911_),
    .X(_00158_));
 sky130_fd_sc_hd__a22o_2 _06594_ (.A1(\tag_array.tag1[13][12] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[14][12] ),
    .X(_03912_));
 sky130_fd_sc_hd__a221o_2 _06595_ (.A1(\tag_array.tag1[12][12] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[15][12] ),
    .C1(_03912_),
    .X(_03913_));
 sky130_fd_sc_hd__a22o_2 _06596_ (.A1(\tag_array.tag1[5][12] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[6][12] ),
    .X(_03914_));
 sky130_fd_sc_hd__a221o_2 _06597_ (.A1(\tag_array.tag1[4][12] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[7][12] ),
    .C1(_03914_),
    .X(_03915_));
 sky130_fd_sc_hd__a22o_2 _06598_ (.A1(\tag_array.tag1[9][12] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[10][12] ),
    .X(_03916_));
 sky130_fd_sc_hd__a221o_2 _06599_ (.A1(\tag_array.tag1[8][12] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[11][12] ),
    .C1(_03916_),
    .X(_03917_));
 sky130_fd_sc_hd__a22o_2 _06600_ (.A1(\tag_array.tag1[1][12] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[2][12] ),
    .X(_03918_));
 sky130_fd_sc_hd__a221o_2 _06601_ (.A1(\tag_array.tag1[0][12] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[3][12] ),
    .C1(_03918_),
    .X(_03919_));
 sky130_fd_sc_hd__a22o_2 _06602_ (.A1(_03522_),
    .A2(_03913_),
    .B1(_03917_),
    .B2(_03506_),
    .X(_03920_));
 sky130_fd_sc_hd__a22o_2 _06603_ (.A1(_03526_),
    .A2(_03915_),
    .B1(_03919_),
    .B2(_03518_),
    .X(_03921_));
 sky130_fd_sc_hd__or2_2 _06604_ (.A(_03920_),
    .B(_03921_),
    .X(_00159_));
 sky130_fd_sc_hd__a22o_2 _06605_ (.A1(\tag_array.tag1[13][13] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[14][13] ),
    .X(_03922_));
 sky130_fd_sc_hd__a221o_2 _06606_ (.A1(\tag_array.tag1[12][13] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[15][13] ),
    .C1(_03922_),
    .X(_03923_));
 sky130_fd_sc_hd__a22o_2 _06607_ (.A1(\tag_array.tag1[5][13] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[6][13] ),
    .X(_03924_));
 sky130_fd_sc_hd__a221o_2 _06608_ (.A1(\tag_array.tag1[4][13] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[7][13] ),
    .C1(_03924_),
    .X(_03925_));
 sky130_fd_sc_hd__a22o_2 _06609_ (.A1(\tag_array.tag1[9][13] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[10][13] ),
    .X(_03926_));
 sky130_fd_sc_hd__a221o_2 _06610_ (.A1(\tag_array.tag1[8][13] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[11][13] ),
    .C1(_03926_),
    .X(_03927_));
 sky130_fd_sc_hd__a22o_2 _06611_ (.A1(\tag_array.tag1[1][13] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[2][13] ),
    .X(_03928_));
 sky130_fd_sc_hd__a221o_2 _06612_ (.A1(\tag_array.tag1[0][13] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[3][13] ),
    .C1(_03928_),
    .X(_03929_));
 sky130_fd_sc_hd__a22o_2 _06613_ (.A1(_03522_),
    .A2(_03923_),
    .B1(_03927_),
    .B2(_03506_),
    .X(_03930_));
 sky130_fd_sc_hd__a22o_2 _06614_ (.A1(_03526_),
    .A2(_03925_),
    .B1(_03929_),
    .B2(_03518_),
    .X(_03931_));
 sky130_fd_sc_hd__or2_2 _06615_ (.A(_03930_),
    .B(_03931_),
    .X(_00160_));
 sky130_fd_sc_hd__a22o_2 _06616_ (.A1(\tag_array.tag1[9][14] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[10][14] ),
    .X(_03932_));
 sky130_fd_sc_hd__a221o_2 _06617_ (.A1(\tag_array.tag1[8][14] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[11][14] ),
    .C1(_03932_),
    .X(_03933_));
 sky130_fd_sc_hd__a22o_2 _06618_ (.A1(\tag_array.tag1[1][14] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[2][14] ),
    .X(_03934_));
 sky130_fd_sc_hd__a221o_2 _06619_ (.A1(\tag_array.tag1[0][14] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[3][14] ),
    .C1(_03934_),
    .X(_03935_));
 sky130_fd_sc_hd__a22o_2 _06620_ (.A1(\tag_array.tag1[13][14] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[14][14] ),
    .X(_03936_));
 sky130_fd_sc_hd__a221o_2 _06621_ (.A1(\tag_array.tag1[12][14] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[15][14] ),
    .C1(_03936_),
    .X(_03937_));
 sky130_fd_sc_hd__a22o_2 _06622_ (.A1(\tag_array.tag1[5][14] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[6][14] ),
    .X(_03938_));
 sky130_fd_sc_hd__a221o_2 _06623_ (.A1(\tag_array.tag1[4][14] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[7][14] ),
    .C1(_03938_),
    .X(_03939_));
 sky130_fd_sc_hd__a22o_2 _06624_ (.A1(_03506_),
    .A2(_03933_),
    .B1(_03937_),
    .B2(_03522_),
    .X(_03940_));
 sky130_fd_sc_hd__a22o_2 _06625_ (.A1(_03518_),
    .A2(_03935_),
    .B1(_03939_),
    .B2(_03526_),
    .X(_03941_));
 sky130_fd_sc_hd__or2_2 _06626_ (.A(_03940_),
    .B(_03941_),
    .X(_00161_));
 sky130_fd_sc_hd__a22o_2 _06627_ (.A1(\tag_array.tag1[9][15] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[10][15] ),
    .X(_03942_));
 sky130_fd_sc_hd__a221o_2 _06628_ (.A1(\tag_array.tag1[8][15] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[11][15] ),
    .C1(_03942_),
    .X(_03943_));
 sky130_fd_sc_hd__a22o_2 _06629_ (.A1(\tag_array.tag1[1][15] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[2][15] ),
    .X(_03944_));
 sky130_fd_sc_hd__a221o_2 _06630_ (.A1(\tag_array.tag1[0][15] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[3][15] ),
    .C1(_03944_),
    .X(_03945_));
 sky130_fd_sc_hd__a22o_2 _06631_ (.A1(\tag_array.tag1[13][15] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[14][15] ),
    .X(_03946_));
 sky130_fd_sc_hd__a221o_2 _06632_ (.A1(\tag_array.tag1[12][15] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[15][15] ),
    .C1(_03946_),
    .X(_03947_));
 sky130_fd_sc_hd__a22o_2 _06633_ (.A1(\tag_array.tag1[5][15] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[6][15] ),
    .X(_03948_));
 sky130_fd_sc_hd__a221o_2 _06634_ (.A1(\tag_array.tag1[4][15] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[7][15] ),
    .C1(_03948_),
    .X(_03949_));
 sky130_fd_sc_hd__a22o_2 _06635_ (.A1(_03506_),
    .A2(_03943_),
    .B1(_03947_),
    .B2(_03522_),
    .X(_03950_));
 sky130_fd_sc_hd__a22o_2 _06636_ (.A1(_03518_),
    .A2(_03945_),
    .B1(_03949_),
    .B2(_03526_),
    .X(_03951_));
 sky130_fd_sc_hd__or2_2 _06637_ (.A(_03950_),
    .B(_03951_),
    .X(_00162_));
 sky130_fd_sc_hd__a22o_2 _06638_ (.A1(\tag_array.tag1[13][16] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[14][16] ),
    .X(_03952_));
 sky130_fd_sc_hd__a221o_2 _06639_ (.A1(\tag_array.tag1[12][16] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[15][16] ),
    .C1(_03952_),
    .X(_03953_));
 sky130_fd_sc_hd__a22o_2 _06640_ (.A1(\tag_array.tag1[1][16] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[2][16] ),
    .X(_03954_));
 sky130_fd_sc_hd__a221o_2 _06641_ (.A1(\tag_array.tag1[0][16] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[3][16] ),
    .C1(_03954_),
    .X(_03955_));
 sky130_fd_sc_hd__a22o_2 _06642_ (.A1(\tag_array.tag1[9][16] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[10][16] ),
    .X(_03956_));
 sky130_fd_sc_hd__a221o_2 _06643_ (.A1(\tag_array.tag1[8][16] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[11][16] ),
    .C1(_03956_),
    .X(_03957_));
 sky130_fd_sc_hd__a22o_2 _06644_ (.A1(\tag_array.tag1[5][16] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[6][16] ),
    .X(_03958_));
 sky130_fd_sc_hd__a221o_2 _06645_ (.A1(\tag_array.tag1[4][16] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[7][16] ),
    .C1(_03958_),
    .X(_03959_));
 sky130_fd_sc_hd__a22o_2 _06646_ (.A1(_03522_),
    .A2(_03953_),
    .B1(_03957_),
    .B2(_03506_),
    .X(_03960_));
 sky130_fd_sc_hd__a22o_2 _06647_ (.A1(_03518_),
    .A2(_03955_),
    .B1(_03959_),
    .B2(_03526_),
    .X(_03961_));
 sky130_fd_sc_hd__or2_2 _06648_ (.A(_03960_),
    .B(_03961_),
    .X(_00163_));
 sky130_fd_sc_hd__a22o_2 _06649_ (.A1(\tag_array.tag1[13][17] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[14][17] ),
    .X(_03962_));
 sky130_fd_sc_hd__a221o_2 _06650_ (.A1(\tag_array.tag1[12][17] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[15][17] ),
    .C1(_03962_),
    .X(_03963_));
 sky130_fd_sc_hd__a22o_2 _06651_ (.A1(\tag_array.tag1[5][17] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[6][17] ),
    .X(_03964_));
 sky130_fd_sc_hd__a221o_2 _06652_ (.A1(\tag_array.tag1[4][17] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[7][17] ),
    .C1(_03964_),
    .X(_03965_));
 sky130_fd_sc_hd__a22o_2 _06653_ (.A1(\tag_array.tag1[9][17] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[10][17] ),
    .X(_03966_));
 sky130_fd_sc_hd__a221o_2 _06654_ (.A1(\tag_array.tag1[8][17] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[11][17] ),
    .C1(_03966_),
    .X(_03967_));
 sky130_fd_sc_hd__a22o_2 _06655_ (.A1(\tag_array.tag1[1][17] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[2][17] ),
    .X(_03968_));
 sky130_fd_sc_hd__a221o_2 _06656_ (.A1(\tag_array.tag1[0][17] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[3][17] ),
    .C1(_03968_),
    .X(_03969_));
 sky130_fd_sc_hd__a22o_2 _06657_ (.A1(_03522_),
    .A2(_03963_),
    .B1(_03967_),
    .B2(_03506_),
    .X(_03970_));
 sky130_fd_sc_hd__a22o_2 _06658_ (.A1(_03526_),
    .A2(_03965_),
    .B1(_03969_),
    .B2(_03518_),
    .X(_03971_));
 sky130_fd_sc_hd__or2_2 _06659_ (.A(_03970_),
    .B(_03971_),
    .X(_00164_));
 sky130_fd_sc_hd__a22o_2 _06660_ (.A1(\tag_array.tag1[13][18] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[14][18] ),
    .X(_03972_));
 sky130_fd_sc_hd__a221o_2 _06661_ (.A1(\tag_array.tag1[12][18] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[15][18] ),
    .C1(_03972_),
    .X(_03973_));
 sky130_fd_sc_hd__a22o_2 _06662_ (.A1(\tag_array.tag1[1][18] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[2][18] ),
    .X(_03974_));
 sky130_fd_sc_hd__a221o_2 _06663_ (.A1(\tag_array.tag1[0][18] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[3][18] ),
    .C1(_03974_),
    .X(_03975_));
 sky130_fd_sc_hd__a22o_2 _06664_ (.A1(\tag_array.tag1[9][18] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[10][18] ),
    .X(_03976_));
 sky130_fd_sc_hd__a221o_2 _06665_ (.A1(\tag_array.tag1[8][18] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[11][18] ),
    .C1(_03976_),
    .X(_03977_));
 sky130_fd_sc_hd__a22o_2 _06666_ (.A1(\tag_array.tag1[5][18] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[6][18] ),
    .X(_03978_));
 sky130_fd_sc_hd__a221o_2 _06667_ (.A1(\tag_array.tag1[4][18] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[7][18] ),
    .C1(_03978_),
    .X(_03979_));
 sky130_fd_sc_hd__a22o_2 _06668_ (.A1(_03522_),
    .A2(_03973_),
    .B1(_03977_),
    .B2(_03506_),
    .X(_03980_));
 sky130_fd_sc_hd__a22o_2 _06669_ (.A1(_03518_),
    .A2(_03975_),
    .B1(_03979_),
    .B2(_03526_),
    .X(_03981_));
 sky130_fd_sc_hd__or2_2 _06670_ (.A(_03980_),
    .B(_03981_),
    .X(_00165_));
 sky130_fd_sc_hd__a22o_2 _06671_ (.A1(\tag_array.tag1[9][19] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[10][19] ),
    .X(_03982_));
 sky130_fd_sc_hd__a221o_2 _06672_ (.A1(\tag_array.tag1[8][19] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[11][19] ),
    .C1(_03982_),
    .X(_03983_));
 sky130_fd_sc_hd__a22o_2 _06673_ (.A1(\tag_array.tag1[5][19] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[6][19] ),
    .X(_03984_));
 sky130_fd_sc_hd__a221o_2 _06674_ (.A1(\tag_array.tag1[4][19] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[7][19] ),
    .C1(_03984_),
    .X(_03985_));
 sky130_fd_sc_hd__a22o_2 _06675_ (.A1(\tag_array.tag1[13][19] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[14][19] ),
    .X(_03986_));
 sky130_fd_sc_hd__a221o_2 _06676_ (.A1(\tag_array.tag1[12][19] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[15][19] ),
    .C1(_03986_),
    .X(_03987_));
 sky130_fd_sc_hd__a22o_2 _06677_ (.A1(\tag_array.tag1[1][19] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[2][19] ),
    .X(_03988_));
 sky130_fd_sc_hd__a221o_2 _06678_ (.A1(\tag_array.tag1[0][19] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[3][19] ),
    .C1(_03988_),
    .X(_03989_));
 sky130_fd_sc_hd__a22o_2 _06679_ (.A1(_03506_),
    .A2(_03983_),
    .B1(_03987_),
    .B2(_03522_),
    .X(_03990_));
 sky130_fd_sc_hd__a22o_2 _06680_ (.A1(_03526_),
    .A2(_03985_),
    .B1(_03989_),
    .B2(_03518_),
    .X(_03991_));
 sky130_fd_sc_hd__or2_2 _06681_ (.A(_03990_),
    .B(_03991_),
    .X(_00166_));
 sky130_fd_sc_hd__a22o_2 _06682_ (.A1(\tag_array.tag1[9][20] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[10][20] ),
    .X(_03992_));
 sky130_fd_sc_hd__a221o_2 _06683_ (.A1(\tag_array.tag1[8][20] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[11][20] ),
    .C1(_03992_),
    .X(_03993_));
 sky130_fd_sc_hd__a22o_2 _06684_ (.A1(\tag_array.tag1[1][20] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[2][20] ),
    .X(_03994_));
 sky130_fd_sc_hd__a221o_2 _06685_ (.A1(\tag_array.tag1[0][20] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[3][20] ),
    .C1(_03994_),
    .X(_03995_));
 sky130_fd_sc_hd__a22o_2 _06686_ (.A1(\tag_array.tag1[13][20] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[14][20] ),
    .X(_03996_));
 sky130_fd_sc_hd__a221o_2 _06687_ (.A1(\tag_array.tag1[12][20] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[15][20] ),
    .C1(_03996_),
    .X(_03997_));
 sky130_fd_sc_hd__a22o_2 _06688_ (.A1(\tag_array.tag1[5][20] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[6][20] ),
    .X(_03998_));
 sky130_fd_sc_hd__a221o_2 _06689_ (.A1(\tag_array.tag1[4][20] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[7][20] ),
    .C1(_03998_),
    .X(_03999_));
 sky130_fd_sc_hd__a22o_2 _06690_ (.A1(_03506_),
    .A2(_03993_),
    .B1(_03997_),
    .B2(_03522_),
    .X(_04000_));
 sky130_fd_sc_hd__a22o_2 _06691_ (.A1(_03518_),
    .A2(_03995_),
    .B1(_03999_),
    .B2(_03526_),
    .X(_04001_));
 sky130_fd_sc_hd__or2_2 _06692_ (.A(_04000_),
    .B(_04001_),
    .X(_00168_));
 sky130_fd_sc_hd__a22o_2 _06693_ (.A1(\tag_array.tag1[9][21] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[10][21] ),
    .X(_04002_));
 sky130_fd_sc_hd__a221o_2 _06694_ (.A1(\tag_array.tag1[8][21] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[11][21] ),
    .C1(_04002_),
    .X(_04003_));
 sky130_fd_sc_hd__a22o_2 _06695_ (.A1(\tag_array.tag1[5][21] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[6][21] ),
    .X(_04004_));
 sky130_fd_sc_hd__a221o_2 _06696_ (.A1(\tag_array.tag1[4][21] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[7][21] ),
    .C1(_04004_),
    .X(_04005_));
 sky130_fd_sc_hd__a22o_2 _06697_ (.A1(\tag_array.tag1[13][21] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[14][21] ),
    .X(_04006_));
 sky130_fd_sc_hd__a221o_2 _06698_ (.A1(\tag_array.tag1[12][21] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[15][21] ),
    .C1(_04006_),
    .X(_04007_));
 sky130_fd_sc_hd__a22o_2 _06699_ (.A1(\tag_array.tag1[1][21] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[2][21] ),
    .X(_04008_));
 sky130_fd_sc_hd__a221o_2 _06700_ (.A1(\tag_array.tag1[0][21] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[3][21] ),
    .C1(_04008_),
    .X(_04009_));
 sky130_fd_sc_hd__a22o_2 _06701_ (.A1(_03506_),
    .A2(_04003_),
    .B1(_04007_),
    .B2(_03522_),
    .X(_04010_));
 sky130_fd_sc_hd__a22o_2 _06702_ (.A1(_03526_),
    .A2(_04005_),
    .B1(_04009_),
    .B2(_03518_),
    .X(_04011_));
 sky130_fd_sc_hd__or2_2 _06703_ (.A(_04010_),
    .B(_04011_),
    .X(_00169_));
 sky130_fd_sc_hd__a22o_2 _06704_ (.A1(\tag_array.tag1[13][22] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[14][22] ),
    .X(_04012_));
 sky130_fd_sc_hd__a221o_2 _06705_ (.A1(\tag_array.tag1[12][22] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[15][22] ),
    .C1(_04012_),
    .X(_04013_));
 sky130_fd_sc_hd__a22o_2 _06706_ (.A1(\tag_array.tag1[1][22] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[2][22] ),
    .X(_04014_));
 sky130_fd_sc_hd__a221o_2 _06707_ (.A1(\tag_array.tag1[0][22] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[3][22] ),
    .C1(_04014_),
    .X(_04015_));
 sky130_fd_sc_hd__a22o_2 _06708_ (.A1(\tag_array.tag1[9][22] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[10][22] ),
    .X(_04016_));
 sky130_fd_sc_hd__a221o_2 _06709_ (.A1(\tag_array.tag1[8][22] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[11][22] ),
    .C1(_04016_),
    .X(_04017_));
 sky130_fd_sc_hd__a22o_2 _06710_ (.A1(\tag_array.tag1[5][22] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[6][22] ),
    .X(_04018_));
 sky130_fd_sc_hd__a221o_2 _06711_ (.A1(\tag_array.tag1[4][22] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[7][22] ),
    .C1(_04018_),
    .X(_04019_));
 sky130_fd_sc_hd__a22o_2 _06712_ (.A1(_03522_),
    .A2(_04013_),
    .B1(_04017_),
    .B2(_03506_),
    .X(_04020_));
 sky130_fd_sc_hd__a22o_2 _06713_ (.A1(_03518_),
    .A2(_04015_),
    .B1(_04019_),
    .B2(_03526_),
    .X(_04021_));
 sky130_fd_sc_hd__or2_2 _06714_ (.A(_04020_),
    .B(_04021_),
    .X(_00170_));
 sky130_fd_sc_hd__a22o_2 _06715_ (.A1(\tag_array.tag1[9][23] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[10][23] ),
    .X(_04022_));
 sky130_fd_sc_hd__a221o_2 _06716_ (.A1(\tag_array.tag1[8][23] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[11][23] ),
    .C1(_04022_),
    .X(_04023_));
 sky130_fd_sc_hd__a22o_2 _06717_ (.A1(\tag_array.tag1[5][23] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[6][23] ),
    .X(_04024_));
 sky130_fd_sc_hd__a221o_2 _06718_ (.A1(\tag_array.tag1[4][23] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[7][23] ),
    .C1(_04024_),
    .X(_04025_));
 sky130_fd_sc_hd__a22o_2 _06719_ (.A1(\tag_array.tag1[13][23] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[14][23] ),
    .X(_04026_));
 sky130_fd_sc_hd__a221o_2 _06720_ (.A1(\tag_array.tag1[12][23] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[15][23] ),
    .C1(_04026_),
    .X(_04027_));
 sky130_fd_sc_hd__a22o_2 _06721_ (.A1(\tag_array.tag1[1][23] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[2][23] ),
    .X(_04028_));
 sky130_fd_sc_hd__a221o_2 _06722_ (.A1(\tag_array.tag1[0][23] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[3][23] ),
    .C1(_04028_),
    .X(_04029_));
 sky130_fd_sc_hd__a22o_2 _06723_ (.A1(_03506_),
    .A2(_04023_),
    .B1(_04027_),
    .B2(_03522_),
    .X(_04030_));
 sky130_fd_sc_hd__a22o_2 _06724_ (.A1(_03526_),
    .A2(_04025_),
    .B1(_04029_),
    .B2(_03518_),
    .X(_04031_));
 sky130_fd_sc_hd__or2_2 _06725_ (.A(_04030_),
    .B(_04031_),
    .X(_00171_));
 sky130_fd_sc_hd__a22o_2 _06726_ (.A1(\tag_array.tag1[13][24] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[14][24] ),
    .X(_04032_));
 sky130_fd_sc_hd__a221o_2 _06727_ (.A1(\tag_array.tag1[12][24] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[15][24] ),
    .C1(_04032_),
    .X(_04033_));
 sky130_fd_sc_hd__a22o_2 _06728_ (.A1(\tag_array.tag1[5][24] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[6][24] ),
    .X(_04034_));
 sky130_fd_sc_hd__a221o_2 _06729_ (.A1(\tag_array.tag1[4][24] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[7][24] ),
    .C1(_04034_),
    .X(_04035_));
 sky130_fd_sc_hd__a22o_2 _06730_ (.A1(\tag_array.tag1[9][24] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[10][24] ),
    .X(_04036_));
 sky130_fd_sc_hd__a221o_2 _06731_ (.A1(\tag_array.tag1[8][24] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[11][24] ),
    .C1(_04036_),
    .X(_04037_));
 sky130_fd_sc_hd__a22o_2 _06732_ (.A1(\tag_array.tag1[1][24] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.tag1[2][24] ),
    .X(_04038_));
 sky130_fd_sc_hd__a221o_2 _06733_ (.A1(\tag_array.tag1[0][24] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.tag1[3][24] ),
    .C1(_04038_),
    .X(_04039_));
 sky130_fd_sc_hd__a22o_2 _06734_ (.A1(_03522_),
    .A2(_04033_),
    .B1(_04037_),
    .B2(_03506_),
    .X(_04040_));
 sky130_fd_sc_hd__a22o_2 _06735_ (.A1(_03526_),
    .A2(_04035_),
    .B1(_04039_),
    .B2(_03518_),
    .X(_04041_));
 sky130_fd_sc_hd__or2_2 _06736_ (.A(_04040_),
    .B(_04041_),
    .X(_00172_));
 sky130_fd_sc_hd__a22o_2 _06737_ (.A1(\data_array.data0[13][0] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][0] ),
    .X(_04042_));
 sky130_fd_sc_hd__a221o_2 _06738_ (.A1(\data_array.data0[12][0] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][0] ),
    .C1(_04042_),
    .X(_04043_));
 sky130_fd_sc_hd__a22o_2 _06739_ (.A1(\data_array.data0[1][0] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][0] ),
    .X(_04044_));
 sky130_fd_sc_hd__a221o_2 _06740_ (.A1(\data_array.data0[0][0] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][0] ),
    .C1(_04044_),
    .X(_04045_));
 sky130_fd_sc_hd__a22o_2 _06741_ (.A1(\data_array.data0[9][0] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][0] ),
    .X(_04046_));
 sky130_fd_sc_hd__a221o_2 _06742_ (.A1(\data_array.data0[8][0] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][0] ),
    .C1(_04046_),
    .X(_04047_));
 sky130_fd_sc_hd__a22o_2 _06743_ (.A1(\data_array.data0[5][0] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][0] ),
    .X(_04048_));
 sky130_fd_sc_hd__a221o_2 _06744_ (.A1(\data_array.data0[4][0] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][0] ),
    .C1(_04048_),
    .X(_04049_));
 sky130_fd_sc_hd__a22o_2 _06745_ (.A1(_03522_),
    .A2(_04043_),
    .B1(_04047_),
    .B2(_03506_),
    .X(_04050_));
 sky130_fd_sc_hd__a22o_2 _06746_ (.A1(_03518_),
    .A2(_04045_),
    .B1(_04049_),
    .B2(_03526_),
    .X(_04051_));
 sky130_fd_sc_hd__or2_2 _06747_ (.A(_04050_),
    .B(_04051_),
    .X(_00000_));
 sky130_fd_sc_hd__a22o_2 _06748_ (.A1(\data_array.data0[13][1] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][1] ),
    .X(_04052_));
 sky130_fd_sc_hd__a221o_2 _06749_ (.A1(\data_array.data0[12][1] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][1] ),
    .C1(_04052_),
    .X(_04053_));
 sky130_fd_sc_hd__a22o_2 _06750_ (.A1(\data_array.data0[1][1] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][1] ),
    .X(_04054_));
 sky130_fd_sc_hd__a221o_2 _06751_ (.A1(\data_array.data0[0][1] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][1] ),
    .C1(_04054_),
    .X(_04055_));
 sky130_fd_sc_hd__a22o_2 _06752_ (.A1(\data_array.data0[9][1] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][1] ),
    .X(_04056_));
 sky130_fd_sc_hd__a221o_2 _06753_ (.A1(\data_array.data0[8][1] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][1] ),
    .C1(_04056_),
    .X(_04057_));
 sky130_fd_sc_hd__a22o_2 _06754_ (.A1(\data_array.data0[5][1] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][1] ),
    .X(_04058_));
 sky130_fd_sc_hd__a221o_2 _06755_ (.A1(\data_array.data0[4][1] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][1] ),
    .C1(_04058_),
    .X(_04059_));
 sky130_fd_sc_hd__a22o_2 _06756_ (.A1(_03522_),
    .A2(_04053_),
    .B1(_04057_),
    .B2(_03506_),
    .X(_04060_));
 sky130_fd_sc_hd__a22o_2 _06757_ (.A1(_03518_),
    .A2(_04055_),
    .B1(_04059_),
    .B2(_03526_),
    .X(_04061_));
 sky130_fd_sc_hd__or2_2 _06758_ (.A(_04060_),
    .B(_04061_),
    .X(_00011_));
 sky130_fd_sc_hd__a22o_2 _06759_ (.A1(\data_array.data0[13][2] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][2] ),
    .X(_04062_));
 sky130_fd_sc_hd__a221o_2 _06760_ (.A1(\data_array.data0[12][2] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][2] ),
    .C1(_04062_),
    .X(_04063_));
 sky130_fd_sc_hd__a22o_2 _06761_ (.A1(\data_array.data0[5][2] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][2] ),
    .X(_04064_));
 sky130_fd_sc_hd__a221o_2 _06762_ (.A1(\data_array.data0[4][2] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][2] ),
    .C1(_04064_),
    .X(_04065_));
 sky130_fd_sc_hd__a22o_2 _06763_ (.A1(\data_array.data0[9][2] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][2] ),
    .X(_04066_));
 sky130_fd_sc_hd__a221o_2 _06764_ (.A1(\data_array.data0[8][2] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][2] ),
    .C1(_04066_),
    .X(_04067_));
 sky130_fd_sc_hd__a22o_2 _06765_ (.A1(\data_array.data0[1][2] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][2] ),
    .X(_04068_));
 sky130_fd_sc_hd__a221o_2 _06766_ (.A1(\data_array.data0[0][2] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][2] ),
    .C1(_04068_),
    .X(_04069_));
 sky130_fd_sc_hd__a22o_2 _06767_ (.A1(_03522_),
    .A2(_04063_),
    .B1(_04067_),
    .B2(_03506_),
    .X(_04070_));
 sky130_fd_sc_hd__a22o_2 _06768_ (.A1(_03526_),
    .A2(_04065_),
    .B1(_04069_),
    .B2(_03518_),
    .X(_04071_));
 sky130_fd_sc_hd__or2_2 _06769_ (.A(_04070_),
    .B(_04071_),
    .X(_00022_));
 sky130_fd_sc_hd__a22o_2 _06770_ (.A1(\data_array.data0[13][3] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][3] ),
    .X(_04072_));
 sky130_fd_sc_hd__a221o_2 _06771_ (.A1(\data_array.data0[12][3] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][3] ),
    .C1(_04072_),
    .X(_04073_));
 sky130_fd_sc_hd__a22o_2 _06772_ (.A1(\data_array.data0[5][3] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][3] ),
    .X(_04074_));
 sky130_fd_sc_hd__a221o_2 _06773_ (.A1(\data_array.data0[4][3] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][3] ),
    .C1(_04074_),
    .X(_04075_));
 sky130_fd_sc_hd__a22o_2 _06774_ (.A1(\data_array.data0[9][3] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][3] ),
    .X(_04076_));
 sky130_fd_sc_hd__a221o_2 _06775_ (.A1(\data_array.data0[8][3] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][3] ),
    .C1(_04076_),
    .X(_04077_));
 sky130_fd_sc_hd__a22o_2 _06776_ (.A1(\data_array.data0[1][3] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][3] ),
    .X(_04078_));
 sky130_fd_sc_hd__a221o_2 _06777_ (.A1(\data_array.data0[0][3] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][3] ),
    .C1(_04078_),
    .X(_04079_));
 sky130_fd_sc_hd__a22o_2 _06778_ (.A1(_03522_),
    .A2(_04073_),
    .B1(_04077_),
    .B2(_03506_),
    .X(_04080_));
 sky130_fd_sc_hd__a22o_2 _06779_ (.A1(_03526_),
    .A2(_04075_),
    .B1(_04079_),
    .B2(_03518_),
    .X(_04081_));
 sky130_fd_sc_hd__or2_2 _06780_ (.A(_04080_),
    .B(_04081_),
    .X(_00033_));
 sky130_fd_sc_hd__a22o_2 _06781_ (.A1(\data_array.data0[9][4] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][4] ),
    .X(_04082_));
 sky130_fd_sc_hd__a221o_2 _06782_ (.A1(\data_array.data0[8][4] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][4] ),
    .C1(_04082_),
    .X(_04083_));
 sky130_fd_sc_hd__a22o_2 _06783_ (.A1(\data_array.data0[5][4] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][4] ),
    .X(_04084_));
 sky130_fd_sc_hd__a221o_2 _06784_ (.A1(\data_array.data0[4][4] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][4] ),
    .C1(_04084_),
    .X(_04085_));
 sky130_fd_sc_hd__a22o_2 _06785_ (.A1(\data_array.data0[13][4] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][4] ),
    .X(_04086_));
 sky130_fd_sc_hd__a221o_2 _06786_ (.A1(\data_array.data0[12][4] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][4] ),
    .C1(_04086_),
    .X(_04087_));
 sky130_fd_sc_hd__a22o_2 _06787_ (.A1(\data_array.data0[1][4] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][4] ),
    .X(_04088_));
 sky130_fd_sc_hd__a221o_2 _06788_ (.A1(\data_array.data0[0][4] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][4] ),
    .C1(_04088_),
    .X(_04089_));
 sky130_fd_sc_hd__a22o_2 _06789_ (.A1(_03506_),
    .A2(_04083_),
    .B1(_04087_),
    .B2(_03522_),
    .X(_04090_));
 sky130_fd_sc_hd__a22o_2 _06790_ (.A1(_03526_),
    .A2(_04085_),
    .B1(_04089_),
    .B2(_03518_),
    .X(_04091_));
 sky130_fd_sc_hd__or2_2 _06791_ (.A(_04090_),
    .B(_04091_),
    .X(_00044_));
 sky130_fd_sc_hd__a22o_2 _06792_ (.A1(\data_array.data0[9][5] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][5] ),
    .X(_04092_));
 sky130_fd_sc_hd__a221o_2 _06793_ (.A1(\data_array.data0[8][5] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][5] ),
    .C1(_04092_),
    .X(_04093_));
 sky130_fd_sc_hd__a22o_2 _06794_ (.A1(\data_array.data0[1][5] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][5] ),
    .X(_04094_));
 sky130_fd_sc_hd__a221o_2 _06795_ (.A1(\data_array.data0[0][5] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][5] ),
    .C1(_04094_),
    .X(_04095_));
 sky130_fd_sc_hd__a22o_2 _06796_ (.A1(\data_array.data0[13][5] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][5] ),
    .X(_04096_));
 sky130_fd_sc_hd__a221o_2 _06797_ (.A1(\data_array.data0[12][5] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][5] ),
    .C1(_04096_),
    .X(_04097_));
 sky130_fd_sc_hd__a22o_2 _06798_ (.A1(\data_array.data0[5][5] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][5] ),
    .X(_04098_));
 sky130_fd_sc_hd__a221o_2 _06799_ (.A1(\data_array.data0[4][5] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][5] ),
    .C1(_04098_),
    .X(_04099_));
 sky130_fd_sc_hd__a22o_2 _06800_ (.A1(_03506_),
    .A2(_04093_),
    .B1(_04097_),
    .B2(_03522_),
    .X(_04100_));
 sky130_fd_sc_hd__a22o_2 _06801_ (.A1(_03518_),
    .A2(_04095_),
    .B1(_04099_),
    .B2(_03526_),
    .X(_04101_));
 sky130_fd_sc_hd__or2_2 _06802_ (.A(_04100_),
    .B(_04101_),
    .X(_00055_));
 sky130_fd_sc_hd__a22o_2 _06803_ (.A1(\data_array.data0[9][6] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][6] ),
    .X(_04102_));
 sky130_fd_sc_hd__a221o_2 _06804_ (.A1(\data_array.data0[8][6] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][6] ),
    .C1(_04102_),
    .X(_04103_));
 sky130_fd_sc_hd__a22o_2 _06805_ (.A1(\data_array.data0[1][6] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][6] ),
    .X(_04104_));
 sky130_fd_sc_hd__a221o_2 _06806_ (.A1(\data_array.data0[0][6] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][6] ),
    .C1(_04104_),
    .X(_04105_));
 sky130_fd_sc_hd__a22o_2 _06807_ (.A1(\data_array.data0[13][6] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][6] ),
    .X(_04106_));
 sky130_fd_sc_hd__a221o_2 _06808_ (.A1(\data_array.data0[12][6] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][6] ),
    .C1(_04106_),
    .X(_04107_));
 sky130_fd_sc_hd__a22o_2 _06809_ (.A1(\data_array.data0[5][6] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][6] ),
    .X(_04108_));
 sky130_fd_sc_hd__a221o_2 _06810_ (.A1(\data_array.data0[4][6] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][6] ),
    .C1(_04108_),
    .X(_04109_));
 sky130_fd_sc_hd__a22o_2 _06811_ (.A1(_03506_),
    .A2(_04103_),
    .B1(_04107_),
    .B2(_03522_),
    .X(_04110_));
 sky130_fd_sc_hd__a22o_2 _06812_ (.A1(_03518_),
    .A2(_04105_),
    .B1(_04109_),
    .B2(_03526_),
    .X(_04111_));
 sky130_fd_sc_hd__or2_2 _06813_ (.A(_04110_),
    .B(_04111_),
    .X(_00060_));
 sky130_fd_sc_hd__a22o_2 _06814_ (.A1(\data_array.data0[9][7] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][7] ),
    .X(_04112_));
 sky130_fd_sc_hd__a221o_2 _06815_ (.A1(\data_array.data0[8][7] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][7] ),
    .C1(_04112_),
    .X(_04113_));
 sky130_fd_sc_hd__a22o_2 _06816_ (.A1(\data_array.data0[1][7] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][7] ),
    .X(_04114_));
 sky130_fd_sc_hd__a221o_2 _06817_ (.A1(\data_array.data0[0][7] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][7] ),
    .C1(_04114_),
    .X(_04115_));
 sky130_fd_sc_hd__a22o_2 _06818_ (.A1(\data_array.data0[13][7] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][7] ),
    .X(_04116_));
 sky130_fd_sc_hd__a221o_2 _06819_ (.A1(\data_array.data0[12][7] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][7] ),
    .C1(_04116_),
    .X(_04117_));
 sky130_fd_sc_hd__a22o_2 _06820_ (.A1(\data_array.data0[5][7] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][7] ),
    .X(_04118_));
 sky130_fd_sc_hd__a221o_2 _06821_ (.A1(\data_array.data0[4][7] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][7] ),
    .C1(_04118_),
    .X(_04119_));
 sky130_fd_sc_hd__a22o_2 _06822_ (.A1(_03506_),
    .A2(_04113_),
    .B1(_04117_),
    .B2(_03522_),
    .X(_04120_));
 sky130_fd_sc_hd__a22o_2 _06823_ (.A1(_03518_),
    .A2(_04115_),
    .B1(_04119_),
    .B2(_03526_),
    .X(_04121_));
 sky130_fd_sc_hd__or2_2 _06824_ (.A(_04120_),
    .B(_04121_),
    .X(_00061_));
 sky130_fd_sc_hd__a22o_2 _06825_ (.A1(\data_array.data0[13][8] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][8] ),
    .X(_04122_));
 sky130_fd_sc_hd__a221o_2 _06826_ (.A1(\data_array.data0[12][8] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][8] ),
    .C1(_04122_),
    .X(_04123_));
 sky130_fd_sc_hd__a22o_2 _06827_ (.A1(\data_array.data0[5][8] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][8] ),
    .X(_04124_));
 sky130_fd_sc_hd__a221o_2 _06828_ (.A1(\data_array.data0[4][8] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][8] ),
    .C1(_04124_),
    .X(_04125_));
 sky130_fd_sc_hd__a22o_2 _06829_ (.A1(\data_array.data0[9][8] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][8] ),
    .X(_04126_));
 sky130_fd_sc_hd__a221o_2 _06830_ (.A1(\data_array.data0[8][8] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][8] ),
    .C1(_04126_),
    .X(_04127_));
 sky130_fd_sc_hd__a22o_2 _06831_ (.A1(\data_array.data0[1][8] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][8] ),
    .X(_04128_));
 sky130_fd_sc_hd__a221o_2 _06832_ (.A1(\data_array.data0[0][8] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][8] ),
    .C1(_04128_),
    .X(_04129_));
 sky130_fd_sc_hd__a22o_2 _06833_ (.A1(_03522_),
    .A2(_04123_),
    .B1(_04127_),
    .B2(_03506_),
    .X(_04130_));
 sky130_fd_sc_hd__a22o_2 _06834_ (.A1(_03526_),
    .A2(_04125_),
    .B1(_04129_),
    .B2(_03518_),
    .X(_04131_));
 sky130_fd_sc_hd__or2_2 _06835_ (.A(_04130_),
    .B(_04131_),
    .X(_00062_));
 sky130_fd_sc_hd__a22o_2 _06836_ (.A1(\data_array.data0[9][9] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][9] ),
    .X(_04132_));
 sky130_fd_sc_hd__a221o_2 _06837_ (.A1(\data_array.data0[8][9] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][9] ),
    .C1(_04132_),
    .X(_04133_));
 sky130_fd_sc_hd__a22o_2 _06838_ (.A1(\data_array.data0[5][9] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][9] ),
    .X(_04134_));
 sky130_fd_sc_hd__a221o_2 _06839_ (.A1(\data_array.data0[4][9] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][9] ),
    .C1(_04134_),
    .X(_04135_));
 sky130_fd_sc_hd__a22o_2 _06840_ (.A1(\data_array.data0[13][9] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][9] ),
    .X(_04136_));
 sky130_fd_sc_hd__a221o_2 _06841_ (.A1(\data_array.data0[12][9] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][9] ),
    .C1(_04136_),
    .X(_04137_));
 sky130_fd_sc_hd__a22o_2 _06842_ (.A1(\data_array.data0[1][9] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][9] ),
    .X(_04138_));
 sky130_fd_sc_hd__a221o_2 _06843_ (.A1(\data_array.data0[0][9] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][9] ),
    .C1(_04138_),
    .X(_04139_));
 sky130_fd_sc_hd__a22o_2 _06844_ (.A1(_03506_),
    .A2(_04133_),
    .B1(_04137_),
    .B2(_03522_),
    .X(_04140_));
 sky130_fd_sc_hd__a22o_2 _06845_ (.A1(_03526_),
    .A2(_04135_),
    .B1(_04139_),
    .B2(_03518_),
    .X(_04141_));
 sky130_fd_sc_hd__or2_2 _06846_ (.A(_04140_),
    .B(_04141_),
    .X(_00063_));
 sky130_fd_sc_hd__a22o_2 _06847_ (.A1(\data_array.data0[9][10] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][10] ),
    .X(_04142_));
 sky130_fd_sc_hd__a221o_2 _06848_ (.A1(\data_array.data0[8][10] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][10] ),
    .C1(_04142_),
    .X(_04143_));
 sky130_fd_sc_hd__a22o_2 _06849_ (.A1(\data_array.data0[5][10] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][10] ),
    .X(_04144_));
 sky130_fd_sc_hd__a221o_2 _06850_ (.A1(\data_array.data0[4][10] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][10] ),
    .C1(_04144_),
    .X(_04145_));
 sky130_fd_sc_hd__a22o_2 _06851_ (.A1(\data_array.data0[13][10] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][10] ),
    .X(_04146_));
 sky130_fd_sc_hd__a221o_2 _06852_ (.A1(\data_array.data0[12][10] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][10] ),
    .C1(_04146_),
    .X(_04147_));
 sky130_fd_sc_hd__a22o_2 _06853_ (.A1(\data_array.data0[1][10] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][10] ),
    .X(_04148_));
 sky130_fd_sc_hd__a221o_2 _06854_ (.A1(\data_array.data0[0][10] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][10] ),
    .C1(_04148_),
    .X(_04149_));
 sky130_fd_sc_hd__a22o_2 _06855_ (.A1(_03506_),
    .A2(_04143_),
    .B1(_04147_),
    .B2(_03522_),
    .X(_04150_));
 sky130_fd_sc_hd__a22o_2 _06856_ (.A1(_03526_),
    .A2(_04145_),
    .B1(_04149_),
    .B2(_03518_),
    .X(_04151_));
 sky130_fd_sc_hd__or2_2 _06857_ (.A(_04150_),
    .B(_04151_),
    .X(_00001_));
 sky130_fd_sc_hd__a22o_2 _06858_ (.A1(\data_array.data0[9][11] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][11] ),
    .X(_04152_));
 sky130_fd_sc_hd__a221o_2 _06859_ (.A1(\data_array.data0[8][11] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][11] ),
    .C1(_04152_),
    .X(_04153_));
 sky130_fd_sc_hd__a22o_2 _06860_ (.A1(\data_array.data0[1][11] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][11] ),
    .X(_04154_));
 sky130_fd_sc_hd__a221o_2 _06861_ (.A1(\data_array.data0[0][11] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][11] ),
    .C1(_04154_),
    .X(_04155_));
 sky130_fd_sc_hd__a22o_2 _06862_ (.A1(\data_array.data0[13][11] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][11] ),
    .X(_04156_));
 sky130_fd_sc_hd__a221o_2 _06863_ (.A1(\data_array.data0[12][11] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][11] ),
    .C1(_04156_),
    .X(_04157_));
 sky130_fd_sc_hd__a22o_2 _06864_ (.A1(\data_array.data0[5][11] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][11] ),
    .X(_04158_));
 sky130_fd_sc_hd__a221o_2 _06865_ (.A1(\data_array.data0[4][11] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][11] ),
    .C1(_04158_),
    .X(_04159_));
 sky130_fd_sc_hd__a22o_2 _06866_ (.A1(_03506_),
    .A2(_04153_),
    .B1(_04157_),
    .B2(_03522_),
    .X(_04160_));
 sky130_fd_sc_hd__a22o_2 _06867_ (.A1(_03518_),
    .A2(_04155_),
    .B1(_04159_),
    .B2(_03526_),
    .X(_04161_));
 sky130_fd_sc_hd__or2_2 _06868_ (.A(_04160_),
    .B(_04161_),
    .X(_00002_));
 sky130_fd_sc_hd__a22o_2 _06869_ (.A1(\data_array.data0[9][12] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][12] ),
    .X(_04162_));
 sky130_fd_sc_hd__a221o_2 _06870_ (.A1(\data_array.data0[8][12] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][12] ),
    .C1(_04162_),
    .X(_04163_));
 sky130_fd_sc_hd__a22o_2 _06871_ (.A1(\data_array.data0[1][12] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][12] ),
    .X(_04164_));
 sky130_fd_sc_hd__a221o_2 _06872_ (.A1(\data_array.data0[0][12] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][12] ),
    .C1(_04164_),
    .X(_04165_));
 sky130_fd_sc_hd__a22o_2 _06873_ (.A1(\data_array.data0[13][12] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][12] ),
    .X(_04166_));
 sky130_fd_sc_hd__a221o_2 _06874_ (.A1(\data_array.data0[12][12] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][12] ),
    .C1(_04166_),
    .X(_04167_));
 sky130_fd_sc_hd__a22o_2 _06875_ (.A1(\data_array.data0[5][12] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][12] ),
    .X(_04168_));
 sky130_fd_sc_hd__a221o_2 _06876_ (.A1(\data_array.data0[4][12] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][12] ),
    .C1(_04168_),
    .X(_04169_));
 sky130_fd_sc_hd__a22o_2 _06877_ (.A1(_03506_),
    .A2(_04163_),
    .B1(_04167_),
    .B2(_03522_),
    .X(_04170_));
 sky130_fd_sc_hd__a22o_2 _06878_ (.A1(_03518_),
    .A2(_04165_),
    .B1(_04169_),
    .B2(_03526_),
    .X(_04171_));
 sky130_fd_sc_hd__or2_2 _06879_ (.A(_04170_),
    .B(_04171_),
    .X(_00003_));
 sky130_fd_sc_hd__a22o_2 _06880_ (.A1(\data_array.data0[13][13] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][13] ),
    .X(_04172_));
 sky130_fd_sc_hd__a221o_2 _06881_ (.A1(\data_array.data0[12][13] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][13] ),
    .C1(_04172_),
    .X(_04173_));
 sky130_fd_sc_hd__a22o_2 _06882_ (.A1(\data_array.data0[1][13] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][13] ),
    .X(_04174_));
 sky130_fd_sc_hd__a221o_2 _06883_ (.A1(\data_array.data0[0][13] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][13] ),
    .C1(_04174_),
    .X(_04175_));
 sky130_fd_sc_hd__a22o_2 _06884_ (.A1(\data_array.data0[9][13] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][13] ),
    .X(_04176_));
 sky130_fd_sc_hd__a221o_2 _06885_ (.A1(\data_array.data0[8][13] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][13] ),
    .C1(_04176_),
    .X(_04177_));
 sky130_fd_sc_hd__a22o_2 _06886_ (.A1(\data_array.data0[5][13] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][13] ),
    .X(_04178_));
 sky130_fd_sc_hd__a221o_2 _06887_ (.A1(\data_array.data0[4][13] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][13] ),
    .C1(_04178_),
    .X(_04179_));
 sky130_fd_sc_hd__a22o_2 _06888_ (.A1(_03522_),
    .A2(_04173_),
    .B1(_04177_),
    .B2(_03506_),
    .X(_04180_));
 sky130_fd_sc_hd__a22o_2 _06889_ (.A1(_03518_),
    .A2(_04175_),
    .B1(_04179_),
    .B2(_03526_),
    .X(_04181_));
 sky130_fd_sc_hd__or2_2 _06890_ (.A(_04180_),
    .B(_04181_),
    .X(_00004_));
 sky130_fd_sc_hd__a22o_2 _06891_ (.A1(\data_array.data0[9][14] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][14] ),
    .X(_04182_));
 sky130_fd_sc_hd__a221o_2 _06892_ (.A1(\data_array.data0[8][14] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][14] ),
    .C1(_04182_),
    .X(_04183_));
 sky130_fd_sc_hd__a22o_2 _06893_ (.A1(\data_array.data0[5][14] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][14] ),
    .X(_04184_));
 sky130_fd_sc_hd__a221o_2 _06894_ (.A1(\data_array.data0[4][14] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][14] ),
    .C1(_04184_),
    .X(_04185_));
 sky130_fd_sc_hd__a22o_2 _06895_ (.A1(\data_array.data0[13][14] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][14] ),
    .X(_04186_));
 sky130_fd_sc_hd__a221o_2 _06896_ (.A1(\data_array.data0[12][14] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][14] ),
    .C1(_04186_),
    .X(_04187_));
 sky130_fd_sc_hd__a22o_2 _06897_ (.A1(\data_array.data0[1][14] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][14] ),
    .X(_04188_));
 sky130_fd_sc_hd__a221o_2 _06898_ (.A1(\data_array.data0[0][14] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][14] ),
    .C1(_04188_),
    .X(_04189_));
 sky130_fd_sc_hd__a22o_2 _06899_ (.A1(_03506_),
    .A2(_04183_),
    .B1(_04187_),
    .B2(_03522_),
    .X(_04190_));
 sky130_fd_sc_hd__a22o_2 _06900_ (.A1(_03526_),
    .A2(_04185_),
    .B1(_04189_),
    .B2(_03518_),
    .X(_04191_));
 sky130_fd_sc_hd__or2_2 _06901_ (.A(_04190_),
    .B(_04191_),
    .X(_00005_));
 sky130_fd_sc_hd__a22o_2 _06902_ (.A1(\data_array.data0[9][15] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][15] ),
    .X(_04192_));
 sky130_fd_sc_hd__a221o_2 _06903_ (.A1(\data_array.data0[8][15] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][15] ),
    .C1(_04192_),
    .X(_04193_));
 sky130_fd_sc_hd__a22o_2 _06904_ (.A1(\data_array.data0[5][15] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][15] ),
    .X(_04194_));
 sky130_fd_sc_hd__a221o_2 _06905_ (.A1(\data_array.data0[4][15] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][15] ),
    .C1(_04194_),
    .X(_04195_));
 sky130_fd_sc_hd__a22o_2 _06906_ (.A1(\data_array.data0[13][15] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][15] ),
    .X(_04196_));
 sky130_fd_sc_hd__a221o_2 _06907_ (.A1(\data_array.data0[12][15] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][15] ),
    .C1(_04196_),
    .X(_04197_));
 sky130_fd_sc_hd__a22o_2 _06908_ (.A1(\data_array.data0[1][15] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][15] ),
    .X(_04198_));
 sky130_fd_sc_hd__a221o_2 _06909_ (.A1(\data_array.data0[0][15] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][15] ),
    .C1(_04198_),
    .X(_04199_));
 sky130_fd_sc_hd__a22o_2 _06910_ (.A1(_03506_),
    .A2(_04193_),
    .B1(_04197_),
    .B2(_03522_),
    .X(_04200_));
 sky130_fd_sc_hd__a22o_2 _06911_ (.A1(_03526_),
    .A2(_04195_),
    .B1(_04199_),
    .B2(_03518_),
    .X(_04201_));
 sky130_fd_sc_hd__or2_2 _06912_ (.A(_04200_),
    .B(_04201_),
    .X(_00006_));
 sky130_fd_sc_hd__a22o_2 _06913_ (.A1(\data_array.data0[9][16] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][16] ),
    .X(_04202_));
 sky130_fd_sc_hd__a221o_2 _06914_ (.A1(\data_array.data0[8][16] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][16] ),
    .C1(_04202_),
    .X(_04203_));
 sky130_fd_sc_hd__a22o_2 _06915_ (.A1(\data_array.data0[5][16] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][16] ),
    .X(_04204_));
 sky130_fd_sc_hd__a221o_2 _06916_ (.A1(\data_array.data0[4][16] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][16] ),
    .C1(_04204_),
    .X(_04205_));
 sky130_fd_sc_hd__a22o_2 _06917_ (.A1(\data_array.data0[13][16] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][16] ),
    .X(_04206_));
 sky130_fd_sc_hd__a221o_2 _06918_ (.A1(\data_array.data0[12][16] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][16] ),
    .C1(_04206_),
    .X(_04207_));
 sky130_fd_sc_hd__a22o_2 _06919_ (.A1(\data_array.data0[1][16] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][16] ),
    .X(_04208_));
 sky130_fd_sc_hd__a221o_2 _06920_ (.A1(\data_array.data0[0][16] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][16] ),
    .C1(_04208_),
    .X(_04209_));
 sky130_fd_sc_hd__a22o_2 _06921_ (.A1(_03506_),
    .A2(_04203_),
    .B1(_04207_),
    .B2(_03522_),
    .X(_04210_));
 sky130_fd_sc_hd__a22o_2 _06922_ (.A1(_03526_),
    .A2(_04205_),
    .B1(_04209_),
    .B2(_03518_),
    .X(_04211_));
 sky130_fd_sc_hd__or2_2 _06923_ (.A(_04210_),
    .B(_04211_),
    .X(_00007_));
 sky130_fd_sc_hd__a22o_2 _06924_ (.A1(\data_array.data0[13][17] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][17] ),
    .X(_04212_));
 sky130_fd_sc_hd__a221o_2 _06925_ (.A1(\data_array.data0[12][17] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][17] ),
    .C1(_04212_),
    .X(_04213_));
 sky130_fd_sc_hd__a22o_2 _06926_ (.A1(\data_array.data0[1][17] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][17] ),
    .X(_04214_));
 sky130_fd_sc_hd__a221o_2 _06927_ (.A1(\data_array.data0[0][17] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][17] ),
    .C1(_04214_),
    .X(_04215_));
 sky130_fd_sc_hd__a22o_2 _06928_ (.A1(\data_array.data0[9][17] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][17] ),
    .X(_04216_));
 sky130_fd_sc_hd__a221o_2 _06929_ (.A1(\data_array.data0[8][17] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][17] ),
    .C1(_04216_),
    .X(_04217_));
 sky130_fd_sc_hd__a22o_2 _06930_ (.A1(\data_array.data0[5][17] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][17] ),
    .X(_04218_));
 sky130_fd_sc_hd__a221o_2 _06931_ (.A1(\data_array.data0[4][17] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][17] ),
    .C1(_04218_),
    .X(_04219_));
 sky130_fd_sc_hd__a22o_2 _06932_ (.A1(_03522_),
    .A2(_04213_),
    .B1(_04217_),
    .B2(_03506_),
    .X(_04220_));
 sky130_fd_sc_hd__a22o_2 _06933_ (.A1(_03518_),
    .A2(_04215_),
    .B1(_04219_),
    .B2(_03526_),
    .X(_04221_));
 sky130_fd_sc_hd__or2_2 _06934_ (.A(_04220_),
    .B(_04221_),
    .X(_00008_));
 sky130_fd_sc_hd__a22o_2 _06935_ (.A1(\data_array.data0[9][18] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][18] ),
    .X(_04222_));
 sky130_fd_sc_hd__a221o_2 _06936_ (.A1(\data_array.data0[8][18] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][18] ),
    .C1(_04222_),
    .X(_04223_));
 sky130_fd_sc_hd__a22o_2 _06937_ (.A1(\data_array.data0[5][18] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][18] ),
    .X(_04224_));
 sky130_fd_sc_hd__a221o_2 _06938_ (.A1(\data_array.data0[4][18] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][18] ),
    .C1(_04224_),
    .X(_04225_));
 sky130_fd_sc_hd__a22o_2 _06939_ (.A1(\data_array.data0[13][18] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][18] ),
    .X(_04226_));
 sky130_fd_sc_hd__a221o_2 _06940_ (.A1(\data_array.data0[12][18] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][18] ),
    .C1(_04226_),
    .X(_04227_));
 sky130_fd_sc_hd__a22o_2 _06941_ (.A1(\data_array.data0[1][18] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][18] ),
    .X(_04228_));
 sky130_fd_sc_hd__a221o_2 _06942_ (.A1(\data_array.data0[0][18] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][18] ),
    .C1(_04228_),
    .X(_04229_));
 sky130_fd_sc_hd__a22o_2 _06943_ (.A1(_03506_),
    .A2(_04223_),
    .B1(_04227_),
    .B2(_03522_),
    .X(_04230_));
 sky130_fd_sc_hd__a22o_2 _06944_ (.A1(_03526_),
    .A2(_04225_),
    .B1(_04229_),
    .B2(_03518_),
    .X(_04231_));
 sky130_fd_sc_hd__or2_2 _06945_ (.A(_04230_),
    .B(_04231_),
    .X(_00009_));
 sky130_fd_sc_hd__a22o_2 _06946_ (.A1(\data_array.data0[13][19] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][19] ),
    .X(_04232_));
 sky130_fd_sc_hd__a221o_2 _06947_ (.A1(\data_array.data0[12][19] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][19] ),
    .C1(_04232_),
    .X(_04233_));
 sky130_fd_sc_hd__a22o_2 _06948_ (.A1(\data_array.data0[5][19] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][19] ),
    .X(_04234_));
 sky130_fd_sc_hd__a221o_2 _06949_ (.A1(\data_array.data0[4][19] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][19] ),
    .C1(_04234_),
    .X(_04235_));
 sky130_fd_sc_hd__a22o_2 _06950_ (.A1(\data_array.data0[9][19] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][19] ),
    .X(_04236_));
 sky130_fd_sc_hd__a221o_2 _06951_ (.A1(\data_array.data0[8][19] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][19] ),
    .C1(_04236_),
    .X(_04237_));
 sky130_fd_sc_hd__a22o_2 _06952_ (.A1(\data_array.data0[1][19] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][19] ),
    .X(_04238_));
 sky130_fd_sc_hd__a221o_2 _06953_ (.A1(\data_array.data0[0][19] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][19] ),
    .C1(_04238_),
    .X(_04239_));
 sky130_fd_sc_hd__a22o_2 _06954_ (.A1(_03522_),
    .A2(_04233_),
    .B1(_04237_),
    .B2(_03506_),
    .X(_04240_));
 sky130_fd_sc_hd__a22o_2 _06955_ (.A1(_03526_),
    .A2(_04235_),
    .B1(_04239_),
    .B2(_03518_),
    .X(_04241_));
 sky130_fd_sc_hd__or2_2 _06956_ (.A(_04240_),
    .B(_04241_),
    .X(_00010_));
 sky130_fd_sc_hd__a22o_2 _06957_ (.A1(\data_array.data0[13][20] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][20] ),
    .X(_04242_));
 sky130_fd_sc_hd__a221o_2 _06958_ (.A1(\data_array.data0[12][20] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][20] ),
    .C1(_04242_),
    .X(_04243_));
 sky130_fd_sc_hd__a22o_2 _06959_ (.A1(\data_array.data0[5][20] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][20] ),
    .X(_04244_));
 sky130_fd_sc_hd__a221o_2 _06960_ (.A1(\data_array.data0[4][20] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][20] ),
    .C1(_04244_),
    .X(_04245_));
 sky130_fd_sc_hd__a22o_2 _06961_ (.A1(\data_array.data0[9][20] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][20] ),
    .X(_04246_));
 sky130_fd_sc_hd__a221o_2 _06962_ (.A1(\data_array.data0[8][20] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][20] ),
    .C1(_04246_),
    .X(_04247_));
 sky130_fd_sc_hd__a22o_2 _06963_ (.A1(\data_array.data0[1][20] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][20] ),
    .X(_04248_));
 sky130_fd_sc_hd__a221o_2 _06964_ (.A1(\data_array.data0[0][20] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][20] ),
    .C1(_04248_),
    .X(_04249_));
 sky130_fd_sc_hd__a22o_2 _06965_ (.A1(_03522_),
    .A2(_04243_),
    .B1(_04247_),
    .B2(_03506_),
    .X(_04250_));
 sky130_fd_sc_hd__a22o_2 _06966_ (.A1(_03526_),
    .A2(_04245_),
    .B1(_04249_),
    .B2(_03518_),
    .X(_04251_));
 sky130_fd_sc_hd__or2_2 _06967_ (.A(_04250_),
    .B(_04251_),
    .X(_00012_));
 sky130_fd_sc_hd__a22o_2 _06968_ (.A1(\data_array.data0[9][21] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][21] ),
    .X(_04252_));
 sky130_fd_sc_hd__a221o_2 _06969_ (.A1(\data_array.data0[8][21] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][21] ),
    .C1(_04252_),
    .X(_04253_));
 sky130_fd_sc_hd__a22o_2 _06970_ (.A1(\data_array.data0[1][21] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][21] ),
    .X(_04254_));
 sky130_fd_sc_hd__a221o_2 _06971_ (.A1(\data_array.data0[0][21] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][21] ),
    .C1(_04254_),
    .X(_04255_));
 sky130_fd_sc_hd__a22o_2 _06972_ (.A1(\data_array.data0[13][21] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][21] ),
    .X(_04256_));
 sky130_fd_sc_hd__a221o_2 _06973_ (.A1(\data_array.data0[12][21] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][21] ),
    .C1(_04256_),
    .X(_04257_));
 sky130_fd_sc_hd__a22o_2 _06974_ (.A1(\data_array.data0[5][21] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][21] ),
    .X(_04258_));
 sky130_fd_sc_hd__a221o_2 _06975_ (.A1(\data_array.data0[4][21] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][21] ),
    .C1(_04258_),
    .X(_04259_));
 sky130_fd_sc_hd__a22o_2 _06976_ (.A1(_03506_),
    .A2(_04253_),
    .B1(_04257_),
    .B2(_03522_),
    .X(_04260_));
 sky130_fd_sc_hd__a22o_2 _06977_ (.A1(_03518_),
    .A2(_04255_),
    .B1(_04259_),
    .B2(_03526_),
    .X(_04261_));
 sky130_fd_sc_hd__or2_2 _06978_ (.A(_04260_),
    .B(_04261_),
    .X(_00013_));
 sky130_fd_sc_hd__a22o_2 _06979_ (.A1(\data_array.data0[9][22] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][22] ),
    .X(_04262_));
 sky130_fd_sc_hd__a221o_2 _06980_ (.A1(\data_array.data0[8][22] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][22] ),
    .C1(_04262_),
    .X(_04263_));
 sky130_fd_sc_hd__a22o_2 _06981_ (.A1(\data_array.data0[1][22] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][22] ),
    .X(_04264_));
 sky130_fd_sc_hd__a221o_2 _06982_ (.A1(\data_array.data0[0][22] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][22] ),
    .C1(_04264_),
    .X(_04265_));
 sky130_fd_sc_hd__a22o_2 _06983_ (.A1(\data_array.data0[13][22] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][22] ),
    .X(_04266_));
 sky130_fd_sc_hd__a221o_2 _06984_ (.A1(\data_array.data0[12][22] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][22] ),
    .C1(_04266_),
    .X(_04267_));
 sky130_fd_sc_hd__a22o_2 _06985_ (.A1(\data_array.data0[5][22] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][22] ),
    .X(_04268_));
 sky130_fd_sc_hd__a221o_2 _06986_ (.A1(\data_array.data0[4][22] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][22] ),
    .C1(_04268_),
    .X(_04269_));
 sky130_fd_sc_hd__a22o_2 _06987_ (.A1(_03506_),
    .A2(_04263_),
    .B1(_04267_),
    .B2(_03522_),
    .X(_04270_));
 sky130_fd_sc_hd__a22o_2 _06988_ (.A1(_03518_),
    .A2(_04265_),
    .B1(_04269_),
    .B2(_03526_),
    .X(_04271_));
 sky130_fd_sc_hd__or2_2 _06989_ (.A(_04270_),
    .B(_04271_),
    .X(_00014_));
 sky130_fd_sc_hd__a22o_2 _06990_ (.A1(\data_array.data0[13][23] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][23] ),
    .X(_04272_));
 sky130_fd_sc_hd__a221o_2 _06991_ (.A1(\data_array.data0[12][23] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][23] ),
    .C1(_04272_),
    .X(_04273_));
 sky130_fd_sc_hd__a22o_2 _06992_ (.A1(\data_array.data0[1][23] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][23] ),
    .X(_04274_));
 sky130_fd_sc_hd__a221o_2 _06993_ (.A1(\data_array.data0[0][23] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][23] ),
    .C1(_04274_),
    .X(_04275_));
 sky130_fd_sc_hd__a22o_2 _06994_ (.A1(\data_array.data0[9][23] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][23] ),
    .X(_04276_));
 sky130_fd_sc_hd__a221o_2 _06995_ (.A1(\data_array.data0[8][23] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][23] ),
    .C1(_04276_),
    .X(_04277_));
 sky130_fd_sc_hd__a22o_2 _06996_ (.A1(\data_array.data0[5][23] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][23] ),
    .X(_04278_));
 sky130_fd_sc_hd__a221o_2 _06997_ (.A1(\data_array.data0[4][23] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][23] ),
    .C1(_04278_),
    .X(_04279_));
 sky130_fd_sc_hd__a22o_2 _06998_ (.A1(_03522_),
    .A2(_04273_),
    .B1(_04277_),
    .B2(_03506_),
    .X(_04280_));
 sky130_fd_sc_hd__a22o_2 _06999_ (.A1(_03518_),
    .A2(_04275_),
    .B1(_04279_),
    .B2(_03526_),
    .X(_04281_));
 sky130_fd_sc_hd__or2_2 _07000_ (.A(_04280_),
    .B(_04281_),
    .X(_00015_));
 sky130_fd_sc_hd__a22o_2 _07001_ (.A1(\data_array.data0[13][24] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][24] ),
    .X(_04282_));
 sky130_fd_sc_hd__a221o_2 _07002_ (.A1(\data_array.data0[12][24] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][24] ),
    .C1(_04282_),
    .X(_04283_));
 sky130_fd_sc_hd__a22o_2 _07003_ (.A1(\data_array.data0[5][24] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][24] ),
    .X(_04284_));
 sky130_fd_sc_hd__a221o_2 _07004_ (.A1(\data_array.data0[4][24] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][24] ),
    .C1(_04284_),
    .X(_04285_));
 sky130_fd_sc_hd__a22o_2 _07005_ (.A1(\data_array.data0[9][24] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][24] ),
    .X(_04286_));
 sky130_fd_sc_hd__a221o_2 _07006_ (.A1(\data_array.data0[8][24] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][24] ),
    .C1(_04286_),
    .X(_04287_));
 sky130_fd_sc_hd__a22o_2 _07007_ (.A1(\data_array.data0[1][24] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][24] ),
    .X(_04288_));
 sky130_fd_sc_hd__a221o_2 _07008_ (.A1(\data_array.data0[0][24] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][24] ),
    .C1(_04288_),
    .X(_04289_));
 sky130_fd_sc_hd__a22o_2 _07009_ (.A1(_03522_),
    .A2(_04283_),
    .B1(_04287_),
    .B2(_03506_),
    .X(_04290_));
 sky130_fd_sc_hd__a22o_2 _07010_ (.A1(_03526_),
    .A2(_04285_),
    .B1(_04289_),
    .B2(_03518_),
    .X(_04291_));
 sky130_fd_sc_hd__or2_2 _07011_ (.A(_04290_),
    .B(_04291_),
    .X(_00016_));
 sky130_fd_sc_hd__a22o_2 _07012_ (.A1(\data_array.data0[13][25] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][25] ),
    .X(_04292_));
 sky130_fd_sc_hd__a221o_2 _07013_ (.A1(\data_array.data0[12][25] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][25] ),
    .C1(_04292_),
    .X(_04293_));
 sky130_fd_sc_hd__a22o_2 _07014_ (.A1(\data_array.data0[1][25] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][25] ),
    .X(_04294_));
 sky130_fd_sc_hd__a221o_2 _07015_ (.A1(\data_array.data0[0][25] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][25] ),
    .C1(_04294_),
    .X(_04295_));
 sky130_fd_sc_hd__a22o_2 _07016_ (.A1(\data_array.data0[9][25] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][25] ),
    .X(_04296_));
 sky130_fd_sc_hd__a221o_2 _07017_ (.A1(\data_array.data0[8][25] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][25] ),
    .C1(_04296_),
    .X(_04297_));
 sky130_fd_sc_hd__a22o_2 _07018_ (.A1(\data_array.data0[5][25] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][25] ),
    .X(_04298_));
 sky130_fd_sc_hd__a221o_2 _07019_ (.A1(\data_array.data0[4][25] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][25] ),
    .C1(_04298_),
    .X(_04299_));
 sky130_fd_sc_hd__a22o_2 _07020_ (.A1(_03522_),
    .A2(_04293_),
    .B1(_04297_),
    .B2(_03506_),
    .X(_04300_));
 sky130_fd_sc_hd__a22o_2 _07021_ (.A1(_03518_),
    .A2(_04295_),
    .B1(_04299_),
    .B2(_03526_),
    .X(_04301_));
 sky130_fd_sc_hd__or2_2 _07022_ (.A(_04300_),
    .B(_04301_),
    .X(_00017_));
 sky130_fd_sc_hd__a22o_2 _07023_ (.A1(\data_array.data0[9][26] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][26] ),
    .X(_04302_));
 sky130_fd_sc_hd__a221o_2 _07024_ (.A1(\data_array.data0[8][26] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][26] ),
    .C1(_04302_),
    .X(_04303_));
 sky130_fd_sc_hd__a22o_2 _07025_ (.A1(\data_array.data0[5][26] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][26] ),
    .X(_04304_));
 sky130_fd_sc_hd__a221o_2 _07026_ (.A1(\data_array.data0[4][26] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][26] ),
    .C1(_04304_),
    .X(_04305_));
 sky130_fd_sc_hd__a22o_2 _07027_ (.A1(\data_array.data0[13][26] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][26] ),
    .X(_04306_));
 sky130_fd_sc_hd__a221o_2 _07028_ (.A1(\data_array.data0[12][26] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][26] ),
    .C1(_04306_),
    .X(_04307_));
 sky130_fd_sc_hd__a22o_2 _07029_ (.A1(\data_array.data0[1][26] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][26] ),
    .X(_04308_));
 sky130_fd_sc_hd__a221o_2 _07030_ (.A1(\data_array.data0[0][26] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][26] ),
    .C1(_04308_),
    .X(_04309_));
 sky130_fd_sc_hd__a22o_2 _07031_ (.A1(_03506_),
    .A2(_04303_),
    .B1(_04307_),
    .B2(_03522_),
    .X(_04310_));
 sky130_fd_sc_hd__a22o_2 _07032_ (.A1(_03526_),
    .A2(_04305_),
    .B1(_04309_),
    .B2(_03518_),
    .X(_04311_));
 sky130_fd_sc_hd__or2_2 _07033_ (.A(_04310_),
    .B(_04311_),
    .X(_00018_));
 sky130_fd_sc_hd__a22o_2 _07034_ (.A1(\data_array.data0[9][27] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][27] ),
    .X(_04312_));
 sky130_fd_sc_hd__a221o_2 _07035_ (.A1(\data_array.data0[8][27] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][27] ),
    .C1(_04312_),
    .X(_04313_));
 sky130_fd_sc_hd__a22o_2 _07036_ (.A1(\data_array.data0[1][27] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][27] ),
    .X(_04314_));
 sky130_fd_sc_hd__a221o_2 _07037_ (.A1(\data_array.data0[0][27] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][27] ),
    .C1(_04314_),
    .X(_04315_));
 sky130_fd_sc_hd__a22o_2 _07038_ (.A1(\data_array.data0[13][27] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][27] ),
    .X(_04316_));
 sky130_fd_sc_hd__a221o_2 _07039_ (.A1(\data_array.data0[12][27] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][27] ),
    .C1(_04316_),
    .X(_04317_));
 sky130_fd_sc_hd__a22o_2 _07040_ (.A1(\data_array.data0[5][27] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][27] ),
    .X(_04318_));
 sky130_fd_sc_hd__a221o_2 _07041_ (.A1(\data_array.data0[4][27] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][27] ),
    .C1(_04318_),
    .X(_04319_));
 sky130_fd_sc_hd__a22o_2 _07042_ (.A1(_03506_),
    .A2(_04313_),
    .B1(_04317_),
    .B2(_03522_),
    .X(_04320_));
 sky130_fd_sc_hd__a22o_2 _07043_ (.A1(_03518_),
    .A2(_04315_),
    .B1(_04319_),
    .B2(_03526_),
    .X(_04321_));
 sky130_fd_sc_hd__or2_2 _07044_ (.A(_04320_),
    .B(_04321_),
    .X(_00019_));
 sky130_fd_sc_hd__a22o_2 _07045_ (.A1(\data_array.data0[9][28] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][28] ),
    .X(_04322_));
 sky130_fd_sc_hd__a221o_2 _07046_ (.A1(\data_array.data0[8][28] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][28] ),
    .C1(_04322_),
    .X(_04323_));
 sky130_fd_sc_hd__a22o_2 _07047_ (.A1(\data_array.data0[5][28] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][28] ),
    .X(_04324_));
 sky130_fd_sc_hd__a221o_2 _07048_ (.A1(\data_array.data0[4][28] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][28] ),
    .C1(_04324_),
    .X(_04325_));
 sky130_fd_sc_hd__a22o_2 _07049_ (.A1(\data_array.data0[13][28] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][28] ),
    .X(_04326_));
 sky130_fd_sc_hd__a221o_2 _07050_ (.A1(\data_array.data0[12][28] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][28] ),
    .C1(_04326_),
    .X(_04327_));
 sky130_fd_sc_hd__a22o_2 _07051_ (.A1(\data_array.data0[1][28] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][28] ),
    .X(_04328_));
 sky130_fd_sc_hd__a221o_2 _07052_ (.A1(\data_array.data0[0][28] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][28] ),
    .C1(_04328_),
    .X(_04329_));
 sky130_fd_sc_hd__a22o_2 _07053_ (.A1(_03506_),
    .A2(_04323_),
    .B1(_04327_),
    .B2(_03522_),
    .X(_04330_));
 sky130_fd_sc_hd__a22o_2 _07054_ (.A1(_03526_),
    .A2(_04325_),
    .B1(_04329_),
    .B2(_03518_),
    .X(_04331_));
 sky130_fd_sc_hd__or2_2 _07055_ (.A(_04330_),
    .B(_04331_),
    .X(_00020_));
 sky130_fd_sc_hd__a22o_2 _07056_ (.A1(\data_array.data0[13][29] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][29] ),
    .X(_04332_));
 sky130_fd_sc_hd__a221o_2 _07057_ (.A1(\data_array.data0[12][29] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][29] ),
    .C1(_04332_),
    .X(_04333_));
 sky130_fd_sc_hd__a22o_2 _07058_ (.A1(\data_array.data0[1][29] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][29] ),
    .X(_04334_));
 sky130_fd_sc_hd__a221o_2 _07059_ (.A1(\data_array.data0[0][29] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][29] ),
    .C1(_04334_),
    .X(_04335_));
 sky130_fd_sc_hd__a22o_2 _07060_ (.A1(\data_array.data0[9][29] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][29] ),
    .X(_04336_));
 sky130_fd_sc_hd__a221o_2 _07061_ (.A1(\data_array.data0[8][29] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][29] ),
    .C1(_04336_),
    .X(_04337_));
 sky130_fd_sc_hd__a22o_2 _07062_ (.A1(\data_array.data0[5][29] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][29] ),
    .X(_04338_));
 sky130_fd_sc_hd__a221o_2 _07063_ (.A1(\data_array.data0[4][29] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][29] ),
    .C1(_04338_),
    .X(_04339_));
 sky130_fd_sc_hd__a22o_2 _07064_ (.A1(_03522_),
    .A2(_04333_),
    .B1(_04337_),
    .B2(_03506_),
    .X(_04340_));
 sky130_fd_sc_hd__a22o_2 _07065_ (.A1(_03518_),
    .A2(_04335_),
    .B1(_04339_),
    .B2(_03526_),
    .X(_04341_));
 sky130_fd_sc_hd__or2_2 _07066_ (.A(_04340_),
    .B(_04341_),
    .X(_00021_));
 sky130_fd_sc_hd__a22o_2 _07067_ (.A1(\data_array.data0[9][30] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][30] ),
    .X(_04342_));
 sky130_fd_sc_hd__a221o_2 _07068_ (.A1(\data_array.data0[8][30] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][30] ),
    .C1(_04342_),
    .X(_04343_));
 sky130_fd_sc_hd__a22o_2 _07069_ (.A1(\data_array.data0[5][30] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][30] ),
    .X(_04344_));
 sky130_fd_sc_hd__a221o_2 _07070_ (.A1(\data_array.data0[4][30] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][30] ),
    .C1(_04344_),
    .X(_04345_));
 sky130_fd_sc_hd__a22o_2 _07071_ (.A1(\data_array.data0[13][30] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][30] ),
    .X(_04346_));
 sky130_fd_sc_hd__a221o_2 _07072_ (.A1(\data_array.data0[12][30] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][30] ),
    .C1(_04346_),
    .X(_04347_));
 sky130_fd_sc_hd__a22o_2 _07073_ (.A1(\data_array.data0[1][30] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][30] ),
    .X(_04348_));
 sky130_fd_sc_hd__a221o_2 _07074_ (.A1(\data_array.data0[0][30] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][30] ),
    .C1(_04348_),
    .X(_04349_));
 sky130_fd_sc_hd__a22o_2 _07075_ (.A1(_03506_),
    .A2(_04343_),
    .B1(_04347_),
    .B2(_03522_),
    .X(_04350_));
 sky130_fd_sc_hd__a22o_2 _07076_ (.A1(_03526_),
    .A2(_04345_),
    .B1(_04349_),
    .B2(_03518_),
    .X(_04351_));
 sky130_fd_sc_hd__or2_2 _07077_ (.A(_04350_),
    .B(_04351_),
    .X(_00023_));
 sky130_fd_sc_hd__a22o_2 _07078_ (.A1(\data_array.data0[13][31] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][31] ),
    .X(_04352_));
 sky130_fd_sc_hd__a221o_2 _07079_ (.A1(\data_array.data0[12][31] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][31] ),
    .C1(_04352_),
    .X(_04353_));
 sky130_fd_sc_hd__a22o_2 _07080_ (.A1(\data_array.data0[5][31] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][31] ),
    .X(_04354_));
 sky130_fd_sc_hd__a221o_2 _07081_ (.A1(\data_array.data0[4][31] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][31] ),
    .C1(_04354_),
    .X(_04355_));
 sky130_fd_sc_hd__a22o_2 _07082_ (.A1(\data_array.data0[9][31] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][31] ),
    .X(_04356_));
 sky130_fd_sc_hd__a221o_2 _07083_ (.A1(\data_array.data0[8][31] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][31] ),
    .C1(_04356_),
    .X(_04357_));
 sky130_fd_sc_hd__a22o_2 _07084_ (.A1(\data_array.data0[1][31] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][31] ),
    .X(_04358_));
 sky130_fd_sc_hd__a221o_2 _07085_ (.A1(\data_array.data0[0][31] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][31] ),
    .C1(_04358_),
    .X(_04359_));
 sky130_fd_sc_hd__a22o_2 _07086_ (.A1(_03522_),
    .A2(_04353_),
    .B1(_04357_),
    .B2(_03506_),
    .X(_04360_));
 sky130_fd_sc_hd__a22o_2 _07087_ (.A1(_03526_),
    .A2(_04355_),
    .B1(_04359_),
    .B2(_03518_),
    .X(_04361_));
 sky130_fd_sc_hd__or2_2 _07088_ (.A(_04360_),
    .B(_04361_),
    .X(_00024_));
 sky130_fd_sc_hd__a22o_2 _07089_ (.A1(\data_array.data0[13][32] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][32] ),
    .X(_04362_));
 sky130_fd_sc_hd__a221o_2 _07090_ (.A1(\data_array.data0[12][32] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][32] ),
    .C1(_04362_),
    .X(_04363_));
 sky130_fd_sc_hd__a22o_2 _07091_ (.A1(\data_array.data0[1][32] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][32] ),
    .X(_04364_));
 sky130_fd_sc_hd__a221o_2 _07092_ (.A1(\data_array.data0[0][32] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][32] ),
    .C1(_04364_),
    .X(_04365_));
 sky130_fd_sc_hd__a22o_2 _07093_ (.A1(\data_array.data0[9][32] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][32] ),
    .X(_04366_));
 sky130_fd_sc_hd__a221o_2 _07094_ (.A1(\data_array.data0[8][32] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][32] ),
    .C1(_04366_),
    .X(_04367_));
 sky130_fd_sc_hd__a22o_2 _07095_ (.A1(\data_array.data0[5][32] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][32] ),
    .X(_04368_));
 sky130_fd_sc_hd__a221o_2 _07096_ (.A1(\data_array.data0[4][32] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][32] ),
    .C1(_04368_),
    .X(_04369_));
 sky130_fd_sc_hd__a22o_2 _07097_ (.A1(_03522_),
    .A2(_04363_),
    .B1(_04367_),
    .B2(_03506_),
    .X(_04370_));
 sky130_fd_sc_hd__a22o_2 _07098_ (.A1(_03518_),
    .A2(_04365_),
    .B1(_04369_),
    .B2(_03526_),
    .X(_04371_));
 sky130_fd_sc_hd__or2_2 _07099_ (.A(_04370_),
    .B(_04371_),
    .X(_00025_));
 sky130_fd_sc_hd__a22o_2 _07100_ (.A1(\data_array.data0[13][33] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][33] ),
    .X(_04372_));
 sky130_fd_sc_hd__a221o_2 _07101_ (.A1(\data_array.data0[12][33] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][33] ),
    .C1(_04372_),
    .X(_04373_));
 sky130_fd_sc_hd__a22o_2 _07102_ (.A1(\data_array.data0[1][33] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][33] ),
    .X(_04374_));
 sky130_fd_sc_hd__a221o_2 _07103_ (.A1(\data_array.data0[0][33] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][33] ),
    .C1(_04374_),
    .X(_04375_));
 sky130_fd_sc_hd__a22o_2 _07104_ (.A1(\data_array.data0[9][33] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][33] ),
    .X(_04376_));
 sky130_fd_sc_hd__a221o_2 _07105_ (.A1(\data_array.data0[8][33] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][33] ),
    .C1(_04376_),
    .X(_04377_));
 sky130_fd_sc_hd__a22o_2 _07106_ (.A1(\data_array.data0[5][33] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][33] ),
    .X(_04378_));
 sky130_fd_sc_hd__a221o_2 _07107_ (.A1(\data_array.data0[4][33] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][33] ),
    .C1(_04378_),
    .X(_04379_));
 sky130_fd_sc_hd__a22o_2 _07108_ (.A1(_03522_),
    .A2(_04373_),
    .B1(_04377_),
    .B2(_03506_),
    .X(_04380_));
 sky130_fd_sc_hd__a22o_2 _07109_ (.A1(_03518_),
    .A2(_04375_),
    .B1(_04379_),
    .B2(_03526_),
    .X(_04381_));
 sky130_fd_sc_hd__or2_2 _07110_ (.A(_04380_),
    .B(_04381_),
    .X(_00026_));
 sky130_fd_sc_hd__a22o_2 _07111_ (.A1(\data_array.data0[13][34] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][34] ),
    .X(_04382_));
 sky130_fd_sc_hd__a221o_2 _07112_ (.A1(\data_array.data0[12][34] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][34] ),
    .C1(_04382_),
    .X(_04383_));
 sky130_fd_sc_hd__a22o_2 _07113_ (.A1(\data_array.data0[5][34] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][34] ),
    .X(_04384_));
 sky130_fd_sc_hd__a221o_2 _07114_ (.A1(\data_array.data0[4][34] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][34] ),
    .C1(_04384_),
    .X(_04385_));
 sky130_fd_sc_hd__a22o_2 _07115_ (.A1(\data_array.data0[9][34] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][34] ),
    .X(_04386_));
 sky130_fd_sc_hd__a221o_2 _07116_ (.A1(\data_array.data0[8][34] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][34] ),
    .C1(_04386_),
    .X(_04387_));
 sky130_fd_sc_hd__a22o_2 _07117_ (.A1(\data_array.data0[1][34] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][34] ),
    .X(_04388_));
 sky130_fd_sc_hd__a221o_2 _07118_ (.A1(\data_array.data0[0][34] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][34] ),
    .C1(_04388_),
    .X(_04389_));
 sky130_fd_sc_hd__a22o_2 _07119_ (.A1(_03522_),
    .A2(_04383_),
    .B1(_04387_),
    .B2(_03506_),
    .X(_04390_));
 sky130_fd_sc_hd__a22o_2 _07120_ (.A1(_03526_),
    .A2(_04385_),
    .B1(_04389_),
    .B2(_03518_),
    .X(_04391_));
 sky130_fd_sc_hd__or2_2 _07121_ (.A(_04390_),
    .B(_04391_),
    .X(_00027_));
 sky130_fd_sc_hd__a22o_2 _07122_ (.A1(\data_array.data0[13][35] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][35] ),
    .X(_04392_));
 sky130_fd_sc_hd__a221o_2 _07123_ (.A1(\data_array.data0[12][35] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][35] ),
    .C1(_04392_),
    .X(_04393_));
 sky130_fd_sc_hd__a22o_2 _07124_ (.A1(\data_array.data0[5][35] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][35] ),
    .X(_04394_));
 sky130_fd_sc_hd__a221o_2 _07125_ (.A1(\data_array.data0[4][35] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][35] ),
    .C1(_04394_),
    .X(_04395_));
 sky130_fd_sc_hd__a22o_2 _07126_ (.A1(\data_array.data0[9][35] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][35] ),
    .X(_04396_));
 sky130_fd_sc_hd__a221o_2 _07127_ (.A1(\data_array.data0[8][35] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][35] ),
    .C1(_04396_),
    .X(_04397_));
 sky130_fd_sc_hd__a22o_2 _07128_ (.A1(\data_array.data0[1][35] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][35] ),
    .X(_04398_));
 sky130_fd_sc_hd__a221o_2 _07129_ (.A1(\data_array.data0[0][35] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][35] ),
    .C1(_04398_),
    .X(_04399_));
 sky130_fd_sc_hd__a22o_2 _07130_ (.A1(_03522_),
    .A2(_04393_),
    .B1(_04397_),
    .B2(_03506_),
    .X(_04400_));
 sky130_fd_sc_hd__a22o_2 _07131_ (.A1(_03526_),
    .A2(_04395_),
    .B1(_04399_),
    .B2(_03518_),
    .X(_04401_));
 sky130_fd_sc_hd__or2_2 _07132_ (.A(_04400_),
    .B(_04401_),
    .X(_00028_));
 sky130_fd_sc_hd__a22o_2 _07133_ (.A1(\data_array.data0[9][36] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][36] ),
    .X(_04402_));
 sky130_fd_sc_hd__a221o_2 _07134_ (.A1(\data_array.data0[8][36] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][36] ),
    .C1(_04402_),
    .X(_04403_));
 sky130_fd_sc_hd__a22o_2 _07135_ (.A1(\data_array.data0[5][36] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][36] ),
    .X(_04404_));
 sky130_fd_sc_hd__a221o_2 _07136_ (.A1(\data_array.data0[4][36] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][36] ),
    .C1(_04404_),
    .X(_04405_));
 sky130_fd_sc_hd__a22o_2 _07137_ (.A1(\data_array.data0[13][36] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][36] ),
    .X(_04406_));
 sky130_fd_sc_hd__a221o_2 _07138_ (.A1(\data_array.data0[12][36] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][36] ),
    .C1(_04406_),
    .X(_04407_));
 sky130_fd_sc_hd__a22o_2 _07139_ (.A1(\data_array.data0[1][36] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][36] ),
    .X(_04408_));
 sky130_fd_sc_hd__a221o_2 _07140_ (.A1(\data_array.data0[0][36] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][36] ),
    .C1(_04408_),
    .X(_04409_));
 sky130_fd_sc_hd__a22o_2 _07141_ (.A1(_03506_),
    .A2(_04403_),
    .B1(_04407_),
    .B2(_03522_),
    .X(_04410_));
 sky130_fd_sc_hd__a22o_2 _07142_ (.A1(_03526_),
    .A2(_04405_),
    .B1(_04409_),
    .B2(_03518_),
    .X(_04411_));
 sky130_fd_sc_hd__or2_2 _07143_ (.A(_04410_),
    .B(_04411_),
    .X(_00029_));
 sky130_fd_sc_hd__a22o_2 _07144_ (.A1(\data_array.data0[9][37] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][37] ),
    .X(_04412_));
 sky130_fd_sc_hd__a221o_2 _07145_ (.A1(\data_array.data0[8][37] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][37] ),
    .C1(_04412_),
    .X(_04413_));
 sky130_fd_sc_hd__a22o_2 _07146_ (.A1(\data_array.data0[1][37] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][37] ),
    .X(_04414_));
 sky130_fd_sc_hd__a221o_2 _07147_ (.A1(\data_array.data0[0][37] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][37] ),
    .C1(_04414_),
    .X(_04415_));
 sky130_fd_sc_hd__a22o_2 _07148_ (.A1(\data_array.data0[13][37] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][37] ),
    .X(_04416_));
 sky130_fd_sc_hd__a221o_2 _07149_ (.A1(\data_array.data0[12][37] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][37] ),
    .C1(_04416_),
    .X(_04417_));
 sky130_fd_sc_hd__a22o_2 _07150_ (.A1(\data_array.data0[5][37] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][37] ),
    .X(_04418_));
 sky130_fd_sc_hd__a221o_2 _07151_ (.A1(\data_array.data0[4][37] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][37] ),
    .C1(_04418_),
    .X(_04419_));
 sky130_fd_sc_hd__a22o_2 _07152_ (.A1(_03506_),
    .A2(_04413_),
    .B1(_04417_),
    .B2(_03522_),
    .X(_04420_));
 sky130_fd_sc_hd__a22o_2 _07153_ (.A1(_03518_),
    .A2(_04415_),
    .B1(_04419_),
    .B2(_03526_),
    .X(_04421_));
 sky130_fd_sc_hd__or2_2 _07154_ (.A(_04420_),
    .B(_04421_),
    .X(_00030_));
 sky130_fd_sc_hd__a22o_2 _07155_ (.A1(\data_array.data0[9][38] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][38] ),
    .X(_04422_));
 sky130_fd_sc_hd__a221o_2 _07156_ (.A1(\data_array.data0[8][38] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][38] ),
    .C1(_04422_),
    .X(_04423_));
 sky130_fd_sc_hd__a22o_2 _07157_ (.A1(\data_array.data0[1][38] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][38] ),
    .X(_04424_));
 sky130_fd_sc_hd__a221o_2 _07158_ (.A1(\data_array.data0[0][38] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][38] ),
    .C1(_04424_),
    .X(_04425_));
 sky130_fd_sc_hd__a22o_2 _07159_ (.A1(\data_array.data0[13][38] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][38] ),
    .X(_04426_));
 sky130_fd_sc_hd__a221o_2 _07160_ (.A1(\data_array.data0[12][38] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][38] ),
    .C1(_04426_),
    .X(_04427_));
 sky130_fd_sc_hd__a22o_2 _07161_ (.A1(\data_array.data0[5][38] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][38] ),
    .X(_04428_));
 sky130_fd_sc_hd__a221o_2 _07162_ (.A1(\data_array.data0[4][38] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][38] ),
    .C1(_04428_),
    .X(_04429_));
 sky130_fd_sc_hd__a22o_2 _07163_ (.A1(_03506_),
    .A2(_04423_),
    .B1(_04427_),
    .B2(_03522_),
    .X(_04430_));
 sky130_fd_sc_hd__a22o_2 _07164_ (.A1(_03518_),
    .A2(_04425_),
    .B1(_04429_),
    .B2(_03526_),
    .X(_04431_));
 sky130_fd_sc_hd__or2_2 _07165_ (.A(_04430_),
    .B(_04431_),
    .X(_00031_));
 sky130_fd_sc_hd__a22o_2 _07166_ (.A1(\data_array.data0[9][39] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][39] ),
    .X(_04432_));
 sky130_fd_sc_hd__a221o_2 _07167_ (.A1(\data_array.data0[8][39] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][39] ),
    .C1(_04432_),
    .X(_04433_));
 sky130_fd_sc_hd__a22o_2 _07168_ (.A1(\data_array.data0[1][39] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][39] ),
    .X(_04434_));
 sky130_fd_sc_hd__a221o_2 _07169_ (.A1(\data_array.data0[0][39] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][39] ),
    .C1(_04434_),
    .X(_04435_));
 sky130_fd_sc_hd__a22o_2 _07170_ (.A1(\data_array.data0[13][39] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][39] ),
    .X(_04436_));
 sky130_fd_sc_hd__a221o_2 _07171_ (.A1(\data_array.data0[12][39] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][39] ),
    .C1(_04436_),
    .X(_04437_));
 sky130_fd_sc_hd__a22o_2 _07172_ (.A1(\data_array.data0[5][39] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][39] ),
    .X(_04438_));
 sky130_fd_sc_hd__a221o_2 _07173_ (.A1(\data_array.data0[4][39] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][39] ),
    .C1(_04438_),
    .X(_04439_));
 sky130_fd_sc_hd__a22o_2 _07174_ (.A1(_03506_),
    .A2(_04433_),
    .B1(_04437_),
    .B2(_03522_),
    .X(_04440_));
 sky130_fd_sc_hd__a22o_2 _07175_ (.A1(_03518_),
    .A2(_04435_),
    .B1(_04439_),
    .B2(_03526_),
    .X(_04441_));
 sky130_fd_sc_hd__or2_2 _07176_ (.A(_04440_),
    .B(_04441_),
    .X(_00032_));
 sky130_fd_sc_hd__a22o_2 _07177_ (.A1(\data_array.data0[13][40] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][40] ),
    .X(_04442_));
 sky130_fd_sc_hd__a221o_2 _07178_ (.A1(\data_array.data0[12][40] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][40] ),
    .C1(_04442_),
    .X(_04443_));
 sky130_fd_sc_hd__a22o_2 _07179_ (.A1(\data_array.data0[5][40] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][40] ),
    .X(_04444_));
 sky130_fd_sc_hd__a221o_2 _07180_ (.A1(\data_array.data0[4][40] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][40] ),
    .C1(_04444_),
    .X(_04445_));
 sky130_fd_sc_hd__a22o_2 _07181_ (.A1(\data_array.data0[9][40] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][40] ),
    .X(_04446_));
 sky130_fd_sc_hd__a221o_2 _07182_ (.A1(\data_array.data0[8][40] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][40] ),
    .C1(_04446_),
    .X(_04447_));
 sky130_fd_sc_hd__a22o_2 _07183_ (.A1(\data_array.data0[1][40] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][40] ),
    .X(_04448_));
 sky130_fd_sc_hd__a221o_2 _07184_ (.A1(\data_array.data0[0][40] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][40] ),
    .C1(_04448_),
    .X(_04449_));
 sky130_fd_sc_hd__a22o_2 _07185_ (.A1(_03522_),
    .A2(_04443_),
    .B1(_04447_),
    .B2(_03506_),
    .X(_04450_));
 sky130_fd_sc_hd__a22o_2 _07186_ (.A1(_03526_),
    .A2(_04445_),
    .B1(_04449_),
    .B2(_03518_),
    .X(_04451_));
 sky130_fd_sc_hd__or2_2 _07187_ (.A(_04450_),
    .B(_04451_),
    .X(_00034_));
 sky130_fd_sc_hd__a22o_2 _07188_ (.A1(\data_array.data0[9][41] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][41] ),
    .X(_04452_));
 sky130_fd_sc_hd__a221o_2 _07189_ (.A1(\data_array.data0[8][41] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][41] ),
    .C1(_04452_),
    .X(_04453_));
 sky130_fd_sc_hd__a22o_2 _07190_ (.A1(\data_array.data0[5][41] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][41] ),
    .X(_04454_));
 sky130_fd_sc_hd__a221o_2 _07191_ (.A1(\data_array.data0[4][41] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][41] ),
    .C1(_04454_),
    .X(_04455_));
 sky130_fd_sc_hd__a22o_2 _07192_ (.A1(\data_array.data0[13][41] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][41] ),
    .X(_04456_));
 sky130_fd_sc_hd__a221o_2 _07193_ (.A1(\data_array.data0[12][41] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][41] ),
    .C1(_04456_),
    .X(_04457_));
 sky130_fd_sc_hd__a22o_2 _07194_ (.A1(\data_array.data0[1][41] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][41] ),
    .X(_04458_));
 sky130_fd_sc_hd__a221o_2 _07195_ (.A1(\data_array.data0[0][41] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][41] ),
    .C1(_04458_),
    .X(_04459_));
 sky130_fd_sc_hd__a22o_2 _07196_ (.A1(_03506_),
    .A2(_04453_),
    .B1(_04457_),
    .B2(_03522_),
    .X(_04460_));
 sky130_fd_sc_hd__a22o_2 _07197_ (.A1(_03526_),
    .A2(_04455_),
    .B1(_04459_),
    .B2(_03518_),
    .X(_04461_));
 sky130_fd_sc_hd__or2_2 _07198_ (.A(_04460_),
    .B(_04461_),
    .X(_00035_));
 sky130_fd_sc_hd__a22o_2 _07199_ (.A1(\data_array.data0[9][42] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][42] ),
    .X(_04462_));
 sky130_fd_sc_hd__a221o_2 _07200_ (.A1(\data_array.data0[8][42] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][42] ),
    .C1(_04462_),
    .X(_04463_));
 sky130_fd_sc_hd__a22o_2 _07201_ (.A1(\data_array.data0[5][42] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][42] ),
    .X(_04464_));
 sky130_fd_sc_hd__a221o_2 _07202_ (.A1(\data_array.data0[4][42] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][42] ),
    .C1(_04464_),
    .X(_04465_));
 sky130_fd_sc_hd__a22o_2 _07203_ (.A1(\data_array.data0[13][42] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][42] ),
    .X(_04466_));
 sky130_fd_sc_hd__a221o_2 _07204_ (.A1(\data_array.data0[12][42] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][42] ),
    .C1(_04466_),
    .X(_04467_));
 sky130_fd_sc_hd__a22o_2 _07205_ (.A1(\data_array.data0[1][42] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][42] ),
    .X(_04468_));
 sky130_fd_sc_hd__a221o_2 _07206_ (.A1(\data_array.data0[0][42] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][42] ),
    .C1(_04468_),
    .X(_04469_));
 sky130_fd_sc_hd__a22o_2 _07207_ (.A1(_03506_),
    .A2(_04463_),
    .B1(_04467_),
    .B2(_03522_),
    .X(_04470_));
 sky130_fd_sc_hd__a22o_2 _07208_ (.A1(_03526_),
    .A2(_04465_),
    .B1(_04469_),
    .B2(_03518_),
    .X(_04471_));
 sky130_fd_sc_hd__or2_2 _07209_ (.A(_04470_),
    .B(_04471_),
    .X(_00036_));
 sky130_fd_sc_hd__a22o_2 _07210_ (.A1(\data_array.data0[9][43] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][43] ),
    .X(_04472_));
 sky130_fd_sc_hd__a221o_2 _07211_ (.A1(\data_array.data0[8][43] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][43] ),
    .C1(_04472_),
    .X(_04473_));
 sky130_fd_sc_hd__a22o_2 _07212_ (.A1(\data_array.data0[1][43] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][43] ),
    .X(_04474_));
 sky130_fd_sc_hd__a221o_2 _07213_ (.A1(\data_array.data0[0][43] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][43] ),
    .C1(_04474_),
    .X(_04475_));
 sky130_fd_sc_hd__a22o_2 _07214_ (.A1(\data_array.data0[13][43] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][43] ),
    .X(_04476_));
 sky130_fd_sc_hd__a221o_2 _07215_ (.A1(\data_array.data0[12][43] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][43] ),
    .C1(_04476_),
    .X(_04477_));
 sky130_fd_sc_hd__a22o_2 _07216_ (.A1(\data_array.data0[5][43] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][43] ),
    .X(_04478_));
 sky130_fd_sc_hd__a221o_2 _07217_ (.A1(\data_array.data0[4][43] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][43] ),
    .C1(_04478_),
    .X(_04479_));
 sky130_fd_sc_hd__a22o_2 _07218_ (.A1(_03506_),
    .A2(_04473_),
    .B1(_04477_),
    .B2(_03522_),
    .X(_04480_));
 sky130_fd_sc_hd__a22o_2 _07219_ (.A1(_03518_),
    .A2(_04475_),
    .B1(_04479_),
    .B2(_03526_),
    .X(_04481_));
 sky130_fd_sc_hd__or2_2 _07220_ (.A(_04480_),
    .B(_04481_),
    .X(_00037_));
 sky130_fd_sc_hd__a22o_2 _07221_ (.A1(\data_array.data0[9][44] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][44] ),
    .X(_04482_));
 sky130_fd_sc_hd__a221o_2 _07222_ (.A1(\data_array.data0[8][44] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][44] ),
    .C1(_04482_),
    .X(_04483_));
 sky130_fd_sc_hd__a22o_2 _07223_ (.A1(\data_array.data0[1][44] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][44] ),
    .X(_04484_));
 sky130_fd_sc_hd__a221o_2 _07224_ (.A1(\data_array.data0[0][44] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][44] ),
    .C1(_04484_),
    .X(_04485_));
 sky130_fd_sc_hd__a22o_2 _07225_ (.A1(\data_array.data0[13][44] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][44] ),
    .X(_04486_));
 sky130_fd_sc_hd__a221o_2 _07226_ (.A1(\data_array.data0[12][44] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][44] ),
    .C1(_04486_),
    .X(_04487_));
 sky130_fd_sc_hd__a22o_2 _07227_ (.A1(\data_array.data0[5][44] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][44] ),
    .X(_04488_));
 sky130_fd_sc_hd__a221o_2 _07228_ (.A1(\data_array.data0[4][44] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][44] ),
    .C1(_04488_),
    .X(_04489_));
 sky130_fd_sc_hd__a22o_2 _07229_ (.A1(_03506_),
    .A2(_04483_),
    .B1(_04487_),
    .B2(_03522_),
    .X(_04490_));
 sky130_fd_sc_hd__a22o_2 _07230_ (.A1(_03518_),
    .A2(_04485_),
    .B1(_04489_),
    .B2(_03526_),
    .X(_04491_));
 sky130_fd_sc_hd__or2_2 _07231_ (.A(_04490_),
    .B(_04491_),
    .X(_00038_));
 sky130_fd_sc_hd__a22o_2 _07232_ (.A1(\data_array.data0[13][45] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][45] ),
    .X(_04492_));
 sky130_fd_sc_hd__a221o_2 _07233_ (.A1(\data_array.data0[12][45] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][45] ),
    .C1(_04492_),
    .X(_04493_));
 sky130_fd_sc_hd__a22o_2 _07234_ (.A1(\data_array.data0[1][45] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][45] ),
    .X(_04494_));
 sky130_fd_sc_hd__a221o_2 _07235_ (.A1(\data_array.data0[0][45] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][45] ),
    .C1(_04494_),
    .X(_04495_));
 sky130_fd_sc_hd__a22o_2 _07236_ (.A1(\data_array.data0[9][45] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][45] ),
    .X(_04496_));
 sky130_fd_sc_hd__a221o_2 _07237_ (.A1(\data_array.data0[8][45] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][45] ),
    .C1(_04496_),
    .X(_04497_));
 sky130_fd_sc_hd__a22o_2 _07238_ (.A1(\data_array.data0[5][45] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][45] ),
    .X(_04498_));
 sky130_fd_sc_hd__a221o_2 _07239_ (.A1(\data_array.data0[4][45] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][45] ),
    .C1(_04498_),
    .X(_04499_));
 sky130_fd_sc_hd__a22o_2 _07240_ (.A1(_03522_),
    .A2(_04493_),
    .B1(_04497_),
    .B2(_03506_),
    .X(_04500_));
 sky130_fd_sc_hd__a22o_2 _07241_ (.A1(_03518_),
    .A2(_04495_),
    .B1(_04499_),
    .B2(_03526_),
    .X(_04501_));
 sky130_fd_sc_hd__or2_2 _07242_ (.A(_04500_),
    .B(_04501_),
    .X(_00039_));
 sky130_fd_sc_hd__a22o_2 _07243_ (.A1(\data_array.data0[9][46] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][46] ),
    .X(_04502_));
 sky130_fd_sc_hd__a221o_2 _07244_ (.A1(\data_array.data0[8][46] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][46] ),
    .C1(_04502_),
    .X(_04503_));
 sky130_fd_sc_hd__a22o_2 _07245_ (.A1(\data_array.data0[5][46] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][46] ),
    .X(_04504_));
 sky130_fd_sc_hd__a221o_2 _07246_ (.A1(\data_array.data0[4][46] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][46] ),
    .C1(_04504_),
    .X(_04505_));
 sky130_fd_sc_hd__a22o_2 _07247_ (.A1(\data_array.data0[13][46] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][46] ),
    .X(_04506_));
 sky130_fd_sc_hd__a221o_2 _07248_ (.A1(\data_array.data0[12][46] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][46] ),
    .C1(_04506_),
    .X(_04507_));
 sky130_fd_sc_hd__a22o_2 _07249_ (.A1(\data_array.data0[1][46] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][46] ),
    .X(_04508_));
 sky130_fd_sc_hd__a221o_2 _07250_ (.A1(\data_array.data0[0][46] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][46] ),
    .C1(_04508_),
    .X(_04509_));
 sky130_fd_sc_hd__a22o_2 _07251_ (.A1(_03506_),
    .A2(_04503_),
    .B1(_04507_),
    .B2(_03522_),
    .X(_04510_));
 sky130_fd_sc_hd__a22o_2 _07252_ (.A1(_03526_),
    .A2(_04505_),
    .B1(_04509_),
    .B2(_03518_),
    .X(_04511_));
 sky130_fd_sc_hd__or2_2 _07253_ (.A(_04510_),
    .B(_04511_),
    .X(_00040_));
 sky130_fd_sc_hd__a22o_2 _07254_ (.A1(\data_array.data0[9][47] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][47] ),
    .X(_04512_));
 sky130_fd_sc_hd__a221o_2 _07255_ (.A1(\data_array.data0[8][47] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][47] ),
    .C1(_04512_),
    .X(_04513_));
 sky130_fd_sc_hd__a22o_2 _07256_ (.A1(\data_array.data0[5][47] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][47] ),
    .X(_04514_));
 sky130_fd_sc_hd__a221o_2 _07257_ (.A1(\data_array.data0[4][47] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][47] ),
    .C1(_04514_),
    .X(_04515_));
 sky130_fd_sc_hd__a22o_2 _07258_ (.A1(\data_array.data0[13][47] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][47] ),
    .X(_04516_));
 sky130_fd_sc_hd__a221o_2 _07259_ (.A1(\data_array.data0[12][47] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][47] ),
    .C1(_04516_),
    .X(_04517_));
 sky130_fd_sc_hd__a22o_2 _07260_ (.A1(\data_array.data0[1][47] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][47] ),
    .X(_04518_));
 sky130_fd_sc_hd__a221o_2 _07261_ (.A1(\data_array.data0[0][47] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][47] ),
    .C1(_04518_),
    .X(_04519_));
 sky130_fd_sc_hd__a22o_2 _07262_ (.A1(_03506_),
    .A2(_04513_),
    .B1(_04517_),
    .B2(_03522_),
    .X(_04520_));
 sky130_fd_sc_hd__a22o_2 _07263_ (.A1(_03526_),
    .A2(_04515_),
    .B1(_04519_),
    .B2(_03518_),
    .X(_04521_));
 sky130_fd_sc_hd__or2_2 _07264_ (.A(_04520_),
    .B(_04521_),
    .X(_00041_));
 sky130_fd_sc_hd__a22o_2 _07265_ (.A1(\data_array.data0[9][48] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][48] ),
    .X(_04522_));
 sky130_fd_sc_hd__a221o_2 _07266_ (.A1(\data_array.data0[8][48] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][48] ),
    .C1(_04522_),
    .X(_04523_));
 sky130_fd_sc_hd__a22o_2 _07267_ (.A1(\data_array.data0[5][48] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][48] ),
    .X(_04524_));
 sky130_fd_sc_hd__a221o_2 _07268_ (.A1(\data_array.data0[4][48] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][48] ),
    .C1(_04524_),
    .X(_04525_));
 sky130_fd_sc_hd__a22o_2 _07269_ (.A1(\data_array.data0[13][48] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][48] ),
    .X(_04526_));
 sky130_fd_sc_hd__a221o_2 _07270_ (.A1(\data_array.data0[12][48] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][48] ),
    .C1(_04526_),
    .X(_04527_));
 sky130_fd_sc_hd__a22o_2 _07271_ (.A1(\data_array.data0[1][48] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][48] ),
    .X(_04528_));
 sky130_fd_sc_hd__a221o_2 _07272_ (.A1(\data_array.data0[0][48] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][48] ),
    .C1(_04528_),
    .X(_04529_));
 sky130_fd_sc_hd__a22o_2 _07273_ (.A1(_03506_),
    .A2(_04523_),
    .B1(_04527_),
    .B2(_03522_),
    .X(_04530_));
 sky130_fd_sc_hd__a22o_2 _07274_ (.A1(_03526_),
    .A2(_04525_),
    .B1(_04529_),
    .B2(_03518_),
    .X(_04531_));
 sky130_fd_sc_hd__or2_2 _07275_ (.A(_04530_),
    .B(_04531_),
    .X(_00042_));
 sky130_fd_sc_hd__a22o_2 _07276_ (.A1(\data_array.data0[13][49] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][49] ),
    .X(_04532_));
 sky130_fd_sc_hd__a221o_2 _07277_ (.A1(\data_array.data0[12][49] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][49] ),
    .C1(_04532_),
    .X(_04533_));
 sky130_fd_sc_hd__a22o_2 _07278_ (.A1(\data_array.data0[1][49] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][49] ),
    .X(_04534_));
 sky130_fd_sc_hd__a221o_2 _07279_ (.A1(\data_array.data0[0][49] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][49] ),
    .C1(_04534_),
    .X(_04535_));
 sky130_fd_sc_hd__a22o_2 _07280_ (.A1(\data_array.data0[9][49] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][49] ),
    .X(_04536_));
 sky130_fd_sc_hd__a221o_2 _07281_ (.A1(\data_array.data0[8][49] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][49] ),
    .C1(_04536_),
    .X(_04537_));
 sky130_fd_sc_hd__a22o_2 _07282_ (.A1(\data_array.data0[5][49] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][49] ),
    .X(_04538_));
 sky130_fd_sc_hd__a221o_2 _07283_ (.A1(\data_array.data0[4][49] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][49] ),
    .C1(_04538_),
    .X(_04539_));
 sky130_fd_sc_hd__a22o_2 _07284_ (.A1(_03522_),
    .A2(_04533_),
    .B1(_04537_),
    .B2(_03506_),
    .X(_04540_));
 sky130_fd_sc_hd__a22o_2 _07285_ (.A1(_03518_),
    .A2(_04535_),
    .B1(_04539_),
    .B2(_03526_),
    .X(_04541_));
 sky130_fd_sc_hd__or2_2 _07286_ (.A(_04540_),
    .B(_04541_),
    .X(_00043_));
 sky130_fd_sc_hd__a22o_2 _07287_ (.A1(\data_array.data0[9][50] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][50] ),
    .X(_04542_));
 sky130_fd_sc_hd__a221o_2 _07288_ (.A1(\data_array.data0[8][50] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][50] ),
    .C1(_04542_),
    .X(_04543_));
 sky130_fd_sc_hd__a22o_2 _07289_ (.A1(\data_array.data0[5][50] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][50] ),
    .X(_04544_));
 sky130_fd_sc_hd__a221o_2 _07290_ (.A1(\data_array.data0[4][50] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][50] ),
    .C1(_04544_),
    .X(_04545_));
 sky130_fd_sc_hd__a22o_2 _07291_ (.A1(\data_array.data0[13][50] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][50] ),
    .X(_04546_));
 sky130_fd_sc_hd__a221o_2 _07292_ (.A1(\data_array.data0[12][50] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][50] ),
    .C1(_04546_),
    .X(_04547_));
 sky130_fd_sc_hd__a22o_2 _07293_ (.A1(\data_array.data0[1][50] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][50] ),
    .X(_04548_));
 sky130_fd_sc_hd__a221o_2 _07294_ (.A1(\data_array.data0[0][50] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][50] ),
    .C1(_04548_),
    .X(_04549_));
 sky130_fd_sc_hd__a22o_2 _07295_ (.A1(_03506_),
    .A2(_04543_),
    .B1(_04547_),
    .B2(_03522_),
    .X(_04550_));
 sky130_fd_sc_hd__a22o_2 _07296_ (.A1(_03526_),
    .A2(_04545_),
    .B1(_04549_),
    .B2(_03518_),
    .X(_04551_));
 sky130_fd_sc_hd__or2_2 _07297_ (.A(_04550_),
    .B(_04551_),
    .X(_00045_));
 sky130_fd_sc_hd__a22o_2 _07298_ (.A1(\data_array.data0[13][51] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][51] ),
    .X(_04552_));
 sky130_fd_sc_hd__a221o_2 _07299_ (.A1(\data_array.data0[12][51] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][51] ),
    .C1(_04552_),
    .X(_04553_));
 sky130_fd_sc_hd__a22o_2 _07300_ (.A1(\data_array.data0[5][51] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][51] ),
    .X(_04554_));
 sky130_fd_sc_hd__a221o_2 _07301_ (.A1(\data_array.data0[4][51] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][51] ),
    .C1(_04554_),
    .X(_04555_));
 sky130_fd_sc_hd__a22o_2 _07302_ (.A1(\data_array.data0[9][51] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][51] ),
    .X(_04556_));
 sky130_fd_sc_hd__a221o_2 _07303_ (.A1(\data_array.data0[8][51] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][51] ),
    .C1(_04556_),
    .X(_04557_));
 sky130_fd_sc_hd__a22o_2 _07304_ (.A1(\data_array.data0[1][51] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][51] ),
    .X(_04558_));
 sky130_fd_sc_hd__a221o_2 _07305_ (.A1(\data_array.data0[0][51] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][51] ),
    .C1(_04558_),
    .X(_04559_));
 sky130_fd_sc_hd__a22o_2 _07306_ (.A1(_03522_),
    .A2(_04553_),
    .B1(_04557_),
    .B2(_03506_),
    .X(_04560_));
 sky130_fd_sc_hd__a22o_2 _07307_ (.A1(_03526_),
    .A2(_04555_),
    .B1(_04559_),
    .B2(_03518_),
    .X(_04561_));
 sky130_fd_sc_hd__or2_2 _07308_ (.A(_04560_),
    .B(_04561_),
    .X(_00046_));
 sky130_fd_sc_hd__a22o_2 _07309_ (.A1(\data_array.data0[13][52] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][52] ),
    .X(_04562_));
 sky130_fd_sc_hd__a221o_2 _07310_ (.A1(\data_array.data0[12][52] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][52] ),
    .C1(_04562_),
    .X(_04563_));
 sky130_fd_sc_hd__a22o_2 _07311_ (.A1(\data_array.data0[5][52] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][52] ),
    .X(_04564_));
 sky130_fd_sc_hd__a221o_2 _07312_ (.A1(\data_array.data0[4][52] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][52] ),
    .C1(_04564_),
    .X(_04565_));
 sky130_fd_sc_hd__a22o_2 _07313_ (.A1(\data_array.data0[9][52] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][52] ),
    .X(_04566_));
 sky130_fd_sc_hd__a221o_2 _07314_ (.A1(\data_array.data0[8][52] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][52] ),
    .C1(_04566_),
    .X(_04567_));
 sky130_fd_sc_hd__a22o_2 _07315_ (.A1(\data_array.data0[1][52] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][52] ),
    .X(_04568_));
 sky130_fd_sc_hd__a221o_2 _07316_ (.A1(\data_array.data0[0][52] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][52] ),
    .C1(_04568_),
    .X(_04569_));
 sky130_fd_sc_hd__a22o_2 _07317_ (.A1(_03522_),
    .A2(_04563_),
    .B1(_04567_),
    .B2(_03506_),
    .X(_04570_));
 sky130_fd_sc_hd__a22o_2 _07318_ (.A1(_03526_),
    .A2(_04565_),
    .B1(_04569_),
    .B2(_03518_),
    .X(_04571_));
 sky130_fd_sc_hd__or2_2 _07319_ (.A(_04570_),
    .B(_04571_),
    .X(_00047_));
 sky130_fd_sc_hd__a22o_2 _07320_ (.A1(\data_array.data0[9][53] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][53] ),
    .X(_04572_));
 sky130_fd_sc_hd__a221o_2 _07321_ (.A1(\data_array.data0[8][53] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][53] ),
    .C1(_04572_),
    .X(_04573_));
 sky130_fd_sc_hd__a22o_2 _07322_ (.A1(\data_array.data0[1][53] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][53] ),
    .X(_04574_));
 sky130_fd_sc_hd__a221o_2 _07323_ (.A1(\data_array.data0[0][53] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][53] ),
    .C1(_04574_),
    .X(_04575_));
 sky130_fd_sc_hd__a22o_2 _07324_ (.A1(\data_array.data0[13][53] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][53] ),
    .X(_04576_));
 sky130_fd_sc_hd__a221o_2 _07325_ (.A1(\data_array.data0[12][53] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][53] ),
    .C1(_04576_),
    .X(_04577_));
 sky130_fd_sc_hd__a22o_2 _07326_ (.A1(\data_array.data0[5][53] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][53] ),
    .X(_04578_));
 sky130_fd_sc_hd__a221o_2 _07327_ (.A1(\data_array.data0[4][53] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][53] ),
    .C1(_04578_),
    .X(_04579_));
 sky130_fd_sc_hd__a22o_2 _07328_ (.A1(_03506_),
    .A2(_04573_),
    .B1(_04577_),
    .B2(_03522_),
    .X(_04580_));
 sky130_fd_sc_hd__a22o_2 _07329_ (.A1(_03518_),
    .A2(_04575_),
    .B1(_04579_),
    .B2(_03526_),
    .X(_04581_));
 sky130_fd_sc_hd__or2_2 _07330_ (.A(_04580_),
    .B(_04581_),
    .X(_00048_));
 sky130_fd_sc_hd__a22o_2 _07331_ (.A1(\data_array.data0[9][54] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][54] ),
    .X(_04582_));
 sky130_fd_sc_hd__a221o_2 _07332_ (.A1(\data_array.data0[8][54] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][54] ),
    .C1(_04582_),
    .X(_04583_));
 sky130_fd_sc_hd__a22o_2 _07333_ (.A1(\data_array.data0[1][54] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][54] ),
    .X(_04584_));
 sky130_fd_sc_hd__a221o_2 _07334_ (.A1(\data_array.data0[0][54] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][54] ),
    .C1(_04584_),
    .X(_04585_));
 sky130_fd_sc_hd__a22o_2 _07335_ (.A1(\data_array.data0[13][54] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][54] ),
    .X(_04586_));
 sky130_fd_sc_hd__a221o_2 _07336_ (.A1(\data_array.data0[12][54] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][54] ),
    .C1(_04586_),
    .X(_04587_));
 sky130_fd_sc_hd__a22o_2 _07337_ (.A1(\data_array.data0[5][54] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][54] ),
    .X(_04588_));
 sky130_fd_sc_hd__a221o_2 _07338_ (.A1(\data_array.data0[4][54] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][54] ),
    .C1(_04588_),
    .X(_04589_));
 sky130_fd_sc_hd__a22o_2 _07339_ (.A1(_03506_),
    .A2(_04583_),
    .B1(_04587_),
    .B2(_03522_),
    .X(_04590_));
 sky130_fd_sc_hd__a22o_2 _07340_ (.A1(_03518_),
    .A2(_04585_),
    .B1(_04589_),
    .B2(_03526_),
    .X(_04591_));
 sky130_fd_sc_hd__or2_2 _07341_ (.A(_04590_),
    .B(_04591_),
    .X(_00049_));
 sky130_fd_sc_hd__a22o_2 _07342_ (.A1(\data_array.data0[13][55] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][55] ),
    .X(_04592_));
 sky130_fd_sc_hd__a221o_2 _07343_ (.A1(\data_array.data0[12][55] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][55] ),
    .C1(_04592_),
    .X(_04593_));
 sky130_fd_sc_hd__a22o_2 _07344_ (.A1(\data_array.data0[1][55] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][55] ),
    .X(_04594_));
 sky130_fd_sc_hd__a221o_2 _07345_ (.A1(\data_array.data0[0][55] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][55] ),
    .C1(_04594_),
    .X(_04595_));
 sky130_fd_sc_hd__a22o_2 _07346_ (.A1(\data_array.data0[9][55] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][55] ),
    .X(_04596_));
 sky130_fd_sc_hd__a221o_2 _07347_ (.A1(\data_array.data0[8][55] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][55] ),
    .C1(_04596_),
    .X(_04597_));
 sky130_fd_sc_hd__a22o_2 _07348_ (.A1(\data_array.data0[5][55] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][55] ),
    .X(_04598_));
 sky130_fd_sc_hd__a221o_2 _07349_ (.A1(\data_array.data0[4][55] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][55] ),
    .C1(_04598_),
    .X(_04599_));
 sky130_fd_sc_hd__a22o_2 _07350_ (.A1(_03522_),
    .A2(_04593_),
    .B1(_04597_),
    .B2(_03506_),
    .X(_04600_));
 sky130_fd_sc_hd__a22o_2 _07351_ (.A1(_03518_),
    .A2(_04595_),
    .B1(_04599_),
    .B2(_03526_),
    .X(_04601_));
 sky130_fd_sc_hd__or2_2 _07352_ (.A(_04600_),
    .B(_04601_),
    .X(_00050_));
 sky130_fd_sc_hd__a22o_2 _07353_ (.A1(\data_array.data0[13][56] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][56] ),
    .X(_04602_));
 sky130_fd_sc_hd__a221o_2 _07354_ (.A1(\data_array.data0[12][56] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][56] ),
    .C1(_04602_),
    .X(_04603_));
 sky130_fd_sc_hd__a22o_2 _07355_ (.A1(\data_array.data0[5][56] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][56] ),
    .X(_04604_));
 sky130_fd_sc_hd__a221o_2 _07356_ (.A1(\data_array.data0[4][56] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][56] ),
    .C1(_04604_),
    .X(_04605_));
 sky130_fd_sc_hd__a22o_2 _07357_ (.A1(\data_array.data0[9][56] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][56] ),
    .X(_04606_));
 sky130_fd_sc_hd__a221o_2 _07358_ (.A1(\data_array.data0[8][56] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][56] ),
    .C1(_04606_),
    .X(_04607_));
 sky130_fd_sc_hd__a22o_2 _07359_ (.A1(\data_array.data0[1][56] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][56] ),
    .X(_04608_));
 sky130_fd_sc_hd__a221o_2 _07360_ (.A1(\data_array.data0[0][56] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][56] ),
    .C1(_04608_),
    .X(_04609_));
 sky130_fd_sc_hd__a22o_2 _07361_ (.A1(_03522_),
    .A2(_04603_),
    .B1(_04607_),
    .B2(_03506_),
    .X(_04610_));
 sky130_fd_sc_hd__a22o_2 _07362_ (.A1(_03526_),
    .A2(_04605_),
    .B1(_04609_),
    .B2(_03518_),
    .X(_04611_));
 sky130_fd_sc_hd__or2_2 _07363_ (.A(_04610_),
    .B(_04611_),
    .X(_00051_));
 sky130_fd_sc_hd__a22o_2 _07364_ (.A1(\data_array.data0[13][57] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][57] ),
    .X(_04612_));
 sky130_fd_sc_hd__a221o_2 _07365_ (.A1(\data_array.data0[12][57] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][57] ),
    .C1(_04612_),
    .X(_04613_));
 sky130_fd_sc_hd__a22o_2 _07366_ (.A1(\data_array.data0[1][57] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][57] ),
    .X(_04614_));
 sky130_fd_sc_hd__a221o_2 _07367_ (.A1(\data_array.data0[0][57] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][57] ),
    .C1(_04614_),
    .X(_04615_));
 sky130_fd_sc_hd__a22o_2 _07368_ (.A1(\data_array.data0[9][57] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][57] ),
    .X(_04616_));
 sky130_fd_sc_hd__a221o_2 _07369_ (.A1(\data_array.data0[8][57] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][57] ),
    .C1(_04616_),
    .X(_04617_));
 sky130_fd_sc_hd__a22o_2 _07370_ (.A1(\data_array.data0[5][57] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][57] ),
    .X(_04618_));
 sky130_fd_sc_hd__a221o_2 _07371_ (.A1(\data_array.data0[4][57] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][57] ),
    .C1(_04618_),
    .X(_04619_));
 sky130_fd_sc_hd__a22o_2 _07372_ (.A1(_03522_),
    .A2(_04613_),
    .B1(_04617_),
    .B2(_03506_),
    .X(_04620_));
 sky130_fd_sc_hd__a22o_2 _07373_ (.A1(_03518_),
    .A2(_04615_),
    .B1(_04619_),
    .B2(_03526_),
    .X(_04621_));
 sky130_fd_sc_hd__or2_2 _07374_ (.A(_04620_),
    .B(_04621_),
    .X(_00052_));
 sky130_fd_sc_hd__a22o_2 _07375_ (.A1(\data_array.data0[9][58] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][58] ),
    .X(_04622_));
 sky130_fd_sc_hd__a221o_2 _07376_ (.A1(\data_array.data0[8][58] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][58] ),
    .C1(_04622_),
    .X(_04623_));
 sky130_fd_sc_hd__a22o_2 _07377_ (.A1(\data_array.data0[5][58] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][58] ),
    .X(_04624_));
 sky130_fd_sc_hd__a221o_2 _07378_ (.A1(\data_array.data0[4][58] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][58] ),
    .C1(_04624_),
    .X(_04625_));
 sky130_fd_sc_hd__a22o_2 _07379_ (.A1(\data_array.data0[13][58] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][58] ),
    .X(_04626_));
 sky130_fd_sc_hd__a221o_2 _07380_ (.A1(\data_array.data0[12][58] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][58] ),
    .C1(_04626_),
    .X(_04627_));
 sky130_fd_sc_hd__a22o_2 _07381_ (.A1(\data_array.data0[1][58] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][58] ),
    .X(_04628_));
 sky130_fd_sc_hd__a221o_2 _07382_ (.A1(\data_array.data0[0][58] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][58] ),
    .C1(_04628_),
    .X(_04629_));
 sky130_fd_sc_hd__a22o_2 _07383_ (.A1(_03506_),
    .A2(_04623_),
    .B1(_04627_),
    .B2(_03522_),
    .X(_04630_));
 sky130_fd_sc_hd__a22o_2 _07384_ (.A1(_03526_),
    .A2(_04625_),
    .B1(_04629_),
    .B2(_03518_),
    .X(_04631_));
 sky130_fd_sc_hd__or2_2 _07385_ (.A(_04630_),
    .B(_04631_),
    .X(_00053_));
 sky130_fd_sc_hd__a22o_2 _07386_ (.A1(\data_array.data0[9][59] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][59] ),
    .X(_04632_));
 sky130_fd_sc_hd__a221o_2 _07387_ (.A1(\data_array.data0[8][59] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][59] ),
    .C1(_04632_),
    .X(_04633_));
 sky130_fd_sc_hd__a22o_2 _07388_ (.A1(\data_array.data0[1][59] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][59] ),
    .X(_04634_));
 sky130_fd_sc_hd__a221o_2 _07389_ (.A1(\data_array.data0[0][59] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][59] ),
    .C1(_04634_),
    .X(_04635_));
 sky130_fd_sc_hd__a22o_2 _07390_ (.A1(\data_array.data0[13][59] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][59] ),
    .X(_04636_));
 sky130_fd_sc_hd__a221o_2 _07391_ (.A1(\data_array.data0[12][59] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][59] ),
    .C1(_04636_),
    .X(_04637_));
 sky130_fd_sc_hd__a22o_2 _07392_ (.A1(\data_array.data0[5][59] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][59] ),
    .X(_04638_));
 sky130_fd_sc_hd__a221o_2 _07393_ (.A1(\data_array.data0[4][59] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][59] ),
    .C1(_04638_),
    .X(_04639_));
 sky130_fd_sc_hd__a22o_2 _07394_ (.A1(_03506_),
    .A2(_04633_),
    .B1(_04637_),
    .B2(_03522_),
    .X(_04640_));
 sky130_fd_sc_hd__a22o_2 _07395_ (.A1(_03518_),
    .A2(_04635_),
    .B1(_04639_),
    .B2(_03526_),
    .X(_04641_));
 sky130_fd_sc_hd__or2_2 _07396_ (.A(_04640_),
    .B(_04641_),
    .X(_00054_));
 sky130_fd_sc_hd__a22o_2 _07397_ (.A1(\data_array.data0[9][60] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][60] ),
    .X(_04642_));
 sky130_fd_sc_hd__a221o_2 _07398_ (.A1(\data_array.data0[8][60] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][60] ),
    .C1(_04642_),
    .X(_04643_));
 sky130_fd_sc_hd__a22o_2 _07399_ (.A1(\data_array.data0[5][60] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][60] ),
    .X(_04644_));
 sky130_fd_sc_hd__a221o_2 _07400_ (.A1(\data_array.data0[4][60] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][60] ),
    .C1(_04644_),
    .X(_04645_));
 sky130_fd_sc_hd__a22o_2 _07401_ (.A1(\data_array.data0[13][60] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][60] ),
    .X(_04646_));
 sky130_fd_sc_hd__a221o_2 _07402_ (.A1(\data_array.data0[12][60] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][60] ),
    .C1(_04646_),
    .X(_04647_));
 sky130_fd_sc_hd__a22o_2 _07403_ (.A1(\data_array.data0[1][60] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][60] ),
    .X(_04648_));
 sky130_fd_sc_hd__a221o_2 _07404_ (.A1(\data_array.data0[0][60] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][60] ),
    .C1(_04648_),
    .X(_04649_));
 sky130_fd_sc_hd__a22o_2 _07405_ (.A1(_03506_),
    .A2(_04643_),
    .B1(_04647_),
    .B2(_03522_),
    .X(_04650_));
 sky130_fd_sc_hd__a22o_2 _07406_ (.A1(_03526_),
    .A2(_04645_),
    .B1(_04649_),
    .B2(_03518_),
    .X(_04651_));
 sky130_fd_sc_hd__or2_2 _07407_ (.A(_04650_),
    .B(_04651_),
    .X(_00056_));
 sky130_fd_sc_hd__a22o_2 _07408_ (.A1(\data_array.data0[13][61] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][61] ),
    .X(_04652_));
 sky130_fd_sc_hd__a221o_2 _07409_ (.A1(\data_array.data0[12][61] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][61] ),
    .C1(_04652_),
    .X(_04653_));
 sky130_fd_sc_hd__a22o_2 _07410_ (.A1(\data_array.data0[1][61] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][61] ),
    .X(_04654_));
 sky130_fd_sc_hd__a221o_2 _07411_ (.A1(\data_array.data0[0][61] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][61] ),
    .C1(_04654_),
    .X(_04655_));
 sky130_fd_sc_hd__a22o_2 _07412_ (.A1(\data_array.data0[9][61] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][61] ),
    .X(_04656_));
 sky130_fd_sc_hd__a221o_2 _07413_ (.A1(\data_array.data0[8][61] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][61] ),
    .C1(_04656_),
    .X(_04657_));
 sky130_fd_sc_hd__a22o_2 _07414_ (.A1(\data_array.data0[5][61] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][61] ),
    .X(_04658_));
 sky130_fd_sc_hd__a221o_2 _07415_ (.A1(\data_array.data0[4][61] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][61] ),
    .C1(_04658_),
    .X(_04659_));
 sky130_fd_sc_hd__a22o_2 _07416_ (.A1(_03522_),
    .A2(_04653_),
    .B1(_04657_),
    .B2(_03506_),
    .X(_04660_));
 sky130_fd_sc_hd__a22o_2 _07417_ (.A1(_03518_),
    .A2(_04655_),
    .B1(_04659_),
    .B2(_03526_),
    .X(_04661_));
 sky130_fd_sc_hd__or2_2 _07418_ (.A(_04660_),
    .B(_04661_),
    .X(_00057_));
 sky130_fd_sc_hd__a22o_2 _07419_ (.A1(\data_array.data0[9][62] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][62] ),
    .X(_04662_));
 sky130_fd_sc_hd__a221o_2 _07420_ (.A1(\data_array.data0[8][62] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][62] ),
    .C1(_04662_),
    .X(_04663_));
 sky130_fd_sc_hd__a22o_2 _07421_ (.A1(\data_array.data0[5][62] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][62] ),
    .X(_04664_));
 sky130_fd_sc_hd__a221o_2 _07422_ (.A1(\data_array.data0[4][62] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][62] ),
    .C1(_04664_),
    .X(_04665_));
 sky130_fd_sc_hd__a22o_2 _07423_ (.A1(\data_array.data0[13][62] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][62] ),
    .X(_04666_));
 sky130_fd_sc_hd__a221o_2 _07424_ (.A1(\data_array.data0[12][62] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][62] ),
    .C1(_04666_),
    .X(_04667_));
 sky130_fd_sc_hd__a22o_2 _07425_ (.A1(\data_array.data0[1][62] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][62] ),
    .X(_04668_));
 sky130_fd_sc_hd__a221o_2 _07426_ (.A1(\data_array.data0[0][62] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][62] ),
    .C1(_04668_),
    .X(_04669_));
 sky130_fd_sc_hd__a22o_2 _07427_ (.A1(_03506_),
    .A2(_04663_),
    .B1(_04667_),
    .B2(_03522_),
    .X(_04670_));
 sky130_fd_sc_hd__a22o_2 _07428_ (.A1(_03526_),
    .A2(_04665_),
    .B1(_04669_),
    .B2(_03518_),
    .X(_04671_));
 sky130_fd_sc_hd__or2_2 _07429_ (.A(_04670_),
    .B(_04671_),
    .X(_00058_));
 sky130_fd_sc_hd__a22o_2 _07430_ (.A1(\data_array.data0[13][63] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[14][63] ),
    .X(_04672_));
 sky130_fd_sc_hd__a221o_2 _07431_ (.A1(\data_array.data0[12][63] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[15][63] ),
    .C1(_04672_),
    .X(_04673_));
 sky130_fd_sc_hd__a22o_2 _07432_ (.A1(\data_array.data0[5][63] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[6][63] ),
    .X(_04674_));
 sky130_fd_sc_hd__a221o_2 _07433_ (.A1(\data_array.data0[4][63] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[7][63] ),
    .C1(_04674_),
    .X(_04675_));
 sky130_fd_sc_hd__a22o_2 _07434_ (.A1(\data_array.data0[9][63] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[10][63] ),
    .X(_04676_));
 sky130_fd_sc_hd__a221o_2 _07435_ (.A1(\data_array.data0[8][63] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[11][63] ),
    .C1(_04676_),
    .X(_04677_));
 sky130_fd_sc_hd__a22o_2 _07436_ (.A1(\data_array.data0[1][63] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data0[2][63] ),
    .X(_04678_));
 sky130_fd_sc_hd__a221o_2 _07437_ (.A1(\data_array.data0[0][63] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data0[3][63] ),
    .C1(_04678_),
    .X(_04679_));
 sky130_fd_sc_hd__a22o_2 _07438_ (.A1(_03522_),
    .A2(_04673_),
    .B1(_04677_),
    .B2(_03506_),
    .X(_04680_));
 sky130_fd_sc_hd__a22o_2 _07439_ (.A1(_03526_),
    .A2(_04675_),
    .B1(_04679_),
    .B2(_03518_),
    .X(_04681_));
 sky130_fd_sc_hd__or2_2 _07440_ (.A(_04680_),
    .B(_04681_),
    .X(_00059_));
 sky130_fd_sc_hd__a22o_2 _07441_ (.A1(\data_array.data1[13][0] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][0] ),
    .X(_04682_));
 sky130_fd_sc_hd__a221o_2 _07442_ (.A1(\data_array.data1[12][0] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][0] ),
    .C1(_04682_),
    .X(_04683_));
 sky130_fd_sc_hd__a22o_2 _07443_ (.A1(\data_array.data1[1][0] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][0] ),
    .X(_04684_));
 sky130_fd_sc_hd__a221o_2 _07444_ (.A1(\data_array.data1[0][0] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][0] ),
    .C1(_04684_),
    .X(_04685_));
 sky130_fd_sc_hd__a22o_2 _07445_ (.A1(\data_array.data1[9][0] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][0] ),
    .X(_04686_));
 sky130_fd_sc_hd__a221o_2 _07446_ (.A1(\data_array.data1[8][0] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][0] ),
    .C1(_04686_),
    .X(_04687_));
 sky130_fd_sc_hd__a22o_2 _07447_ (.A1(\data_array.data1[5][0] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][0] ),
    .X(_04688_));
 sky130_fd_sc_hd__a221o_2 _07448_ (.A1(\data_array.data1[4][0] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][0] ),
    .C1(_04688_),
    .X(_04689_));
 sky130_fd_sc_hd__a22o_2 _07449_ (.A1(_03522_),
    .A2(_04683_),
    .B1(_04687_),
    .B2(_03506_),
    .X(_04690_));
 sky130_fd_sc_hd__a22o_2 _07450_ (.A1(_03518_),
    .A2(_04685_),
    .B1(_04689_),
    .B2(_03526_),
    .X(_04691_));
 sky130_fd_sc_hd__or2_2 _07451_ (.A(_04690_),
    .B(_04691_),
    .X(_00064_));
 sky130_fd_sc_hd__a22o_2 _07452_ (.A1(\data_array.data1[13][1] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][1] ),
    .X(_04692_));
 sky130_fd_sc_hd__a221o_2 _07453_ (.A1(\data_array.data1[12][1] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][1] ),
    .C1(_04692_),
    .X(_04693_));
 sky130_fd_sc_hd__a22o_2 _07454_ (.A1(\data_array.data1[1][1] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][1] ),
    .X(_04694_));
 sky130_fd_sc_hd__a221o_2 _07455_ (.A1(\data_array.data1[0][1] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][1] ),
    .C1(_04694_),
    .X(_04695_));
 sky130_fd_sc_hd__a22o_2 _07456_ (.A1(\data_array.data1[9][1] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][1] ),
    .X(_04696_));
 sky130_fd_sc_hd__a221o_2 _07457_ (.A1(\data_array.data1[8][1] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][1] ),
    .C1(_04696_),
    .X(_04697_));
 sky130_fd_sc_hd__a22o_2 _07458_ (.A1(\data_array.data1[5][1] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][1] ),
    .X(_04698_));
 sky130_fd_sc_hd__a221o_2 _07459_ (.A1(\data_array.data1[4][1] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][1] ),
    .C1(_04698_),
    .X(_04699_));
 sky130_fd_sc_hd__a22o_2 _07460_ (.A1(_03522_),
    .A2(_04693_),
    .B1(_04697_),
    .B2(_03506_),
    .X(_04700_));
 sky130_fd_sc_hd__a22o_2 _07461_ (.A1(_03518_),
    .A2(_04695_),
    .B1(_04699_),
    .B2(_03526_),
    .X(_04701_));
 sky130_fd_sc_hd__or2_2 _07462_ (.A(_04700_),
    .B(_04701_),
    .X(_00075_));
 sky130_fd_sc_hd__a22o_2 _07463_ (.A1(\data_array.data1[13][2] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][2] ),
    .X(_04702_));
 sky130_fd_sc_hd__a221o_2 _07464_ (.A1(\data_array.data1[12][2] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][2] ),
    .C1(_04702_),
    .X(_04703_));
 sky130_fd_sc_hd__a22o_2 _07465_ (.A1(\data_array.data1[5][2] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][2] ),
    .X(_04704_));
 sky130_fd_sc_hd__a221o_2 _07466_ (.A1(\data_array.data1[4][2] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][2] ),
    .C1(_04704_),
    .X(_04705_));
 sky130_fd_sc_hd__a22o_2 _07467_ (.A1(\data_array.data1[9][2] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][2] ),
    .X(_04706_));
 sky130_fd_sc_hd__a221o_2 _07468_ (.A1(\data_array.data1[8][2] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][2] ),
    .C1(_04706_),
    .X(_04707_));
 sky130_fd_sc_hd__a22o_2 _07469_ (.A1(\data_array.data1[1][2] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][2] ),
    .X(_04708_));
 sky130_fd_sc_hd__a221o_2 _07470_ (.A1(\data_array.data1[0][2] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][2] ),
    .C1(_04708_),
    .X(_04709_));
 sky130_fd_sc_hd__a22o_2 _07471_ (.A1(_03522_),
    .A2(_04703_),
    .B1(_04707_),
    .B2(_03506_),
    .X(_04710_));
 sky130_fd_sc_hd__a22o_2 _07472_ (.A1(_03526_),
    .A2(_04705_),
    .B1(_04709_),
    .B2(_03518_),
    .X(_04711_));
 sky130_fd_sc_hd__or2_2 _07473_ (.A(_04710_),
    .B(_04711_),
    .X(_00086_));
 sky130_fd_sc_hd__a22o_2 _07474_ (.A1(\data_array.data1[13][3] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][3] ),
    .X(_04712_));
 sky130_fd_sc_hd__a221o_2 _07475_ (.A1(\data_array.data1[12][3] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][3] ),
    .C1(_04712_),
    .X(_04713_));
 sky130_fd_sc_hd__a22o_2 _07476_ (.A1(\data_array.data1[5][3] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][3] ),
    .X(_04714_));
 sky130_fd_sc_hd__a221o_2 _07477_ (.A1(\data_array.data1[4][3] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][3] ),
    .C1(_04714_),
    .X(_04715_));
 sky130_fd_sc_hd__a22o_2 _07478_ (.A1(\data_array.data1[9][3] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][3] ),
    .X(_04716_));
 sky130_fd_sc_hd__a221o_2 _07479_ (.A1(\data_array.data1[8][3] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][3] ),
    .C1(_04716_),
    .X(_04717_));
 sky130_fd_sc_hd__a22o_2 _07480_ (.A1(\data_array.data1[1][3] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][3] ),
    .X(_04718_));
 sky130_fd_sc_hd__a221o_2 _07481_ (.A1(\data_array.data1[0][3] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][3] ),
    .C1(_04718_),
    .X(_04719_));
 sky130_fd_sc_hd__a22o_2 _07482_ (.A1(_03522_),
    .A2(_04713_),
    .B1(_04717_),
    .B2(_03506_),
    .X(_04720_));
 sky130_fd_sc_hd__a22o_2 _07483_ (.A1(_03526_),
    .A2(_04715_),
    .B1(_04719_),
    .B2(_03518_),
    .X(_04721_));
 sky130_fd_sc_hd__or2_2 _07484_ (.A(_04720_),
    .B(_04721_),
    .X(_00097_));
 sky130_fd_sc_hd__a22o_2 _07485_ (.A1(\data_array.data1[9][4] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][4] ),
    .X(_04722_));
 sky130_fd_sc_hd__a221o_2 _07486_ (.A1(\data_array.data1[8][4] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][4] ),
    .C1(_04722_),
    .X(_04723_));
 sky130_fd_sc_hd__a22o_2 _07487_ (.A1(\data_array.data1[5][4] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][4] ),
    .X(_04724_));
 sky130_fd_sc_hd__a221o_2 _07488_ (.A1(\data_array.data1[4][4] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][4] ),
    .C1(_04724_),
    .X(_04725_));
 sky130_fd_sc_hd__a22o_2 _07489_ (.A1(\data_array.data1[13][4] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][4] ),
    .X(_04726_));
 sky130_fd_sc_hd__a221o_2 _07490_ (.A1(\data_array.data1[12][4] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][4] ),
    .C1(_04726_),
    .X(_04727_));
 sky130_fd_sc_hd__a22o_2 _07491_ (.A1(\data_array.data1[1][4] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][4] ),
    .X(_04728_));
 sky130_fd_sc_hd__a221o_2 _07492_ (.A1(\data_array.data1[0][4] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][4] ),
    .C1(_04728_),
    .X(_04729_));
 sky130_fd_sc_hd__a22o_2 _07493_ (.A1(_03506_),
    .A2(_04723_),
    .B1(_04727_),
    .B2(_03522_),
    .X(_04730_));
 sky130_fd_sc_hd__a22o_2 _07494_ (.A1(_03526_),
    .A2(_04725_),
    .B1(_04729_),
    .B2(_03518_),
    .X(_04731_));
 sky130_fd_sc_hd__or2_2 _07495_ (.A(_04730_),
    .B(_04731_),
    .X(_00108_));
 sky130_fd_sc_hd__a22o_2 _07496_ (.A1(\data_array.data1[9][5] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][5] ),
    .X(_04732_));
 sky130_fd_sc_hd__a221o_2 _07497_ (.A1(\data_array.data1[8][5] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][5] ),
    .C1(_04732_),
    .X(_04733_));
 sky130_fd_sc_hd__a22o_2 _07498_ (.A1(\data_array.data1[1][5] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][5] ),
    .X(_04734_));
 sky130_fd_sc_hd__a221o_2 _07499_ (.A1(\data_array.data1[0][5] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][5] ),
    .C1(_04734_),
    .X(_04735_));
 sky130_fd_sc_hd__a22o_2 _07500_ (.A1(\data_array.data1[13][5] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][5] ),
    .X(_04736_));
 sky130_fd_sc_hd__a221o_2 _07501_ (.A1(\data_array.data1[12][5] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][5] ),
    .C1(_04736_),
    .X(_04737_));
 sky130_fd_sc_hd__a22o_2 _07502_ (.A1(\data_array.data1[5][5] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][5] ),
    .X(_04738_));
 sky130_fd_sc_hd__a221o_2 _07503_ (.A1(\data_array.data1[4][5] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][5] ),
    .C1(_04738_),
    .X(_04739_));
 sky130_fd_sc_hd__a22o_2 _07504_ (.A1(_03506_),
    .A2(_04733_),
    .B1(_04737_),
    .B2(_03522_),
    .X(_04740_));
 sky130_fd_sc_hd__a22o_2 _07505_ (.A1(_03518_),
    .A2(_04735_),
    .B1(_04739_),
    .B2(_03526_),
    .X(_04741_));
 sky130_fd_sc_hd__or2_2 _07506_ (.A(_04740_),
    .B(_04741_),
    .X(_00119_));
 sky130_fd_sc_hd__a22o_2 _07507_ (.A1(\data_array.data1[9][6] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][6] ),
    .X(_04742_));
 sky130_fd_sc_hd__a221o_2 _07508_ (.A1(\data_array.data1[8][6] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][6] ),
    .C1(_04742_),
    .X(_04743_));
 sky130_fd_sc_hd__a22o_2 _07509_ (.A1(\data_array.data1[1][6] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][6] ),
    .X(_04744_));
 sky130_fd_sc_hd__a221o_2 _07510_ (.A1(\data_array.data1[0][6] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][6] ),
    .C1(_04744_),
    .X(_04745_));
 sky130_fd_sc_hd__a22o_2 _07511_ (.A1(\data_array.data1[13][6] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][6] ),
    .X(_04746_));
 sky130_fd_sc_hd__a221o_2 _07512_ (.A1(\data_array.data1[12][6] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][6] ),
    .C1(_04746_),
    .X(_04747_));
 sky130_fd_sc_hd__a22o_2 _07513_ (.A1(\data_array.data1[5][6] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][6] ),
    .X(_04748_));
 sky130_fd_sc_hd__a221o_2 _07514_ (.A1(\data_array.data1[4][6] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][6] ),
    .C1(_04748_),
    .X(_04749_));
 sky130_fd_sc_hd__a22o_2 _07515_ (.A1(_03506_),
    .A2(_04743_),
    .B1(_04747_),
    .B2(_03522_),
    .X(_04750_));
 sky130_fd_sc_hd__a22o_2 _07516_ (.A1(_03518_),
    .A2(_04745_),
    .B1(_04749_),
    .B2(_03526_),
    .X(_04751_));
 sky130_fd_sc_hd__or2_2 _07517_ (.A(_04750_),
    .B(_04751_),
    .X(_00124_));
 sky130_fd_sc_hd__a22o_2 _07518_ (.A1(\data_array.data1[9][7] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][7] ),
    .X(_04752_));
 sky130_fd_sc_hd__a221o_2 _07519_ (.A1(\data_array.data1[8][7] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][7] ),
    .C1(_04752_),
    .X(_04753_));
 sky130_fd_sc_hd__a22o_2 _07520_ (.A1(\data_array.data1[1][7] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][7] ),
    .X(_04754_));
 sky130_fd_sc_hd__a221o_2 _07521_ (.A1(\data_array.data1[0][7] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][7] ),
    .C1(_04754_),
    .X(_04755_));
 sky130_fd_sc_hd__a22o_2 _07522_ (.A1(\data_array.data1[13][7] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][7] ),
    .X(_04756_));
 sky130_fd_sc_hd__a221o_2 _07523_ (.A1(\data_array.data1[12][7] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][7] ),
    .C1(_04756_),
    .X(_04757_));
 sky130_fd_sc_hd__a22o_2 _07524_ (.A1(\data_array.data1[5][7] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][7] ),
    .X(_04758_));
 sky130_fd_sc_hd__a221o_2 _07525_ (.A1(\data_array.data1[4][7] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][7] ),
    .C1(_04758_),
    .X(_04759_));
 sky130_fd_sc_hd__a22o_2 _07526_ (.A1(_03506_),
    .A2(_04753_),
    .B1(_04757_),
    .B2(_03522_),
    .X(_04760_));
 sky130_fd_sc_hd__a22o_2 _07527_ (.A1(_03518_),
    .A2(_04755_),
    .B1(_04759_),
    .B2(_03526_),
    .X(_04761_));
 sky130_fd_sc_hd__or2_2 _07528_ (.A(_04760_),
    .B(_04761_),
    .X(_00125_));
 sky130_fd_sc_hd__a22o_2 _07529_ (.A1(\data_array.data1[13][8] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][8] ),
    .X(_04762_));
 sky130_fd_sc_hd__a221o_2 _07530_ (.A1(\data_array.data1[12][8] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][8] ),
    .C1(_04762_),
    .X(_04763_));
 sky130_fd_sc_hd__a22o_2 _07531_ (.A1(\data_array.data1[5][8] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][8] ),
    .X(_04764_));
 sky130_fd_sc_hd__a221o_2 _07532_ (.A1(\data_array.data1[4][8] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][8] ),
    .C1(_04764_),
    .X(_04765_));
 sky130_fd_sc_hd__a22o_2 _07533_ (.A1(\data_array.data1[9][8] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][8] ),
    .X(_04766_));
 sky130_fd_sc_hd__a221o_2 _07534_ (.A1(\data_array.data1[8][8] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][8] ),
    .C1(_04766_),
    .X(_04767_));
 sky130_fd_sc_hd__a22o_2 _07535_ (.A1(\data_array.data1[1][8] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][8] ),
    .X(_04768_));
 sky130_fd_sc_hd__a221o_2 _07536_ (.A1(\data_array.data1[0][8] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][8] ),
    .C1(_04768_),
    .X(_04769_));
 sky130_fd_sc_hd__a22o_2 _07537_ (.A1(_03522_),
    .A2(_04763_),
    .B1(_04767_),
    .B2(_03506_),
    .X(_04770_));
 sky130_fd_sc_hd__a22o_2 _07538_ (.A1(_03526_),
    .A2(_04765_),
    .B1(_04769_),
    .B2(_03518_),
    .X(_04771_));
 sky130_fd_sc_hd__or2_2 _07539_ (.A(_04770_),
    .B(_04771_),
    .X(_00126_));
 sky130_fd_sc_hd__a22o_2 _07540_ (.A1(\data_array.data1[9][9] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][9] ),
    .X(_04772_));
 sky130_fd_sc_hd__a221o_2 _07541_ (.A1(\data_array.data1[8][9] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][9] ),
    .C1(_04772_),
    .X(_04773_));
 sky130_fd_sc_hd__a22o_2 _07542_ (.A1(\data_array.data1[5][9] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][9] ),
    .X(_04774_));
 sky130_fd_sc_hd__a221o_2 _07543_ (.A1(\data_array.data1[4][9] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][9] ),
    .C1(_04774_),
    .X(_04775_));
 sky130_fd_sc_hd__a22o_2 _07544_ (.A1(\data_array.data1[13][9] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][9] ),
    .X(_04776_));
 sky130_fd_sc_hd__a221o_2 _07545_ (.A1(\data_array.data1[12][9] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][9] ),
    .C1(_04776_),
    .X(_04777_));
 sky130_fd_sc_hd__a22o_2 _07546_ (.A1(\data_array.data1[1][9] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][9] ),
    .X(_04778_));
 sky130_fd_sc_hd__a221o_2 _07547_ (.A1(\data_array.data1[0][9] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][9] ),
    .C1(_04778_),
    .X(_04779_));
 sky130_fd_sc_hd__a22o_2 _07548_ (.A1(_03506_),
    .A2(_04773_),
    .B1(_04777_),
    .B2(_03522_),
    .X(_04780_));
 sky130_fd_sc_hd__a22o_2 _07549_ (.A1(_03526_),
    .A2(_04775_),
    .B1(_04779_),
    .B2(_03518_),
    .X(_04781_));
 sky130_fd_sc_hd__or2_2 _07550_ (.A(_04780_),
    .B(_04781_),
    .X(_00127_));
 sky130_fd_sc_hd__a22o_2 _07551_ (.A1(\data_array.data1[9][10] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][10] ),
    .X(_04782_));
 sky130_fd_sc_hd__a221o_2 _07552_ (.A1(\data_array.data1[8][10] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][10] ),
    .C1(_04782_),
    .X(_04783_));
 sky130_fd_sc_hd__a22o_2 _07553_ (.A1(\data_array.data1[5][10] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][10] ),
    .X(_04784_));
 sky130_fd_sc_hd__a221o_2 _07554_ (.A1(\data_array.data1[4][10] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][10] ),
    .C1(_04784_),
    .X(_04785_));
 sky130_fd_sc_hd__a22o_2 _07555_ (.A1(\data_array.data1[13][10] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][10] ),
    .X(_04786_));
 sky130_fd_sc_hd__a221o_2 _07556_ (.A1(\data_array.data1[12][10] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][10] ),
    .C1(_04786_),
    .X(_04787_));
 sky130_fd_sc_hd__a22o_2 _07557_ (.A1(\data_array.data1[1][10] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][10] ),
    .X(_04788_));
 sky130_fd_sc_hd__a221o_2 _07558_ (.A1(\data_array.data1[0][10] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][10] ),
    .C1(_04788_),
    .X(_04789_));
 sky130_fd_sc_hd__a22o_2 _07559_ (.A1(_03506_),
    .A2(_04783_),
    .B1(_04787_),
    .B2(_03522_),
    .X(_04790_));
 sky130_fd_sc_hd__a22o_2 _07560_ (.A1(_03526_),
    .A2(_04785_),
    .B1(_04789_),
    .B2(_03518_),
    .X(_04791_));
 sky130_fd_sc_hd__or2_2 _07561_ (.A(_04790_),
    .B(_04791_),
    .X(_00065_));
 sky130_fd_sc_hd__a22o_2 _07562_ (.A1(\data_array.data1[9][11] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][11] ),
    .X(_04792_));
 sky130_fd_sc_hd__a221o_2 _07563_ (.A1(\data_array.data1[8][11] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][11] ),
    .C1(_04792_),
    .X(_04793_));
 sky130_fd_sc_hd__a22o_2 _07564_ (.A1(\data_array.data1[1][11] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][11] ),
    .X(_04794_));
 sky130_fd_sc_hd__a221o_2 _07565_ (.A1(\data_array.data1[0][11] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][11] ),
    .C1(_04794_),
    .X(_04795_));
 sky130_fd_sc_hd__a22o_2 _07566_ (.A1(\data_array.data1[13][11] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][11] ),
    .X(_04796_));
 sky130_fd_sc_hd__a221o_2 _07567_ (.A1(\data_array.data1[12][11] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][11] ),
    .C1(_04796_),
    .X(_04797_));
 sky130_fd_sc_hd__a22o_2 _07568_ (.A1(\data_array.data1[5][11] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][11] ),
    .X(_04798_));
 sky130_fd_sc_hd__a221o_2 _07569_ (.A1(\data_array.data1[4][11] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][11] ),
    .C1(_04798_),
    .X(_04799_));
 sky130_fd_sc_hd__a22o_2 _07570_ (.A1(_03506_),
    .A2(_04793_),
    .B1(_04797_),
    .B2(_03522_),
    .X(_04800_));
 sky130_fd_sc_hd__a22o_2 _07571_ (.A1(_03518_),
    .A2(_04795_),
    .B1(_04799_),
    .B2(_03526_),
    .X(_04801_));
 sky130_fd_sc_hd__or2_2 _07572_ (.A(_04800_),
    .B(_04801_),
    .X(_00066_));
 sky130_fd_sc_hd__a22o_2 _07573_ (.A1(\data_array.data1[9][12] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][12] ),
    .X(_04802_));
 sky130_fd_sc_hd__a221o_2 _07574_ (.A1(\data_array.data1[8][12] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][12] ),
    .C1(_04802_),
    .X(_04803_));
 sky130_fd_sc_hd__a22o_2 _07575_ (.A1(\data_array.data1[1][12] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][12] ),
    .X(_04804_));
 sky130_fd_sc_hd__a221o_2 _07576_ (.A1(\data_array.data1[0][12] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][12] ),
    .C1(_04804_),
    .X(_04805_));
 sky130_fd_sc_hd__a22o_2 _07577_ (.A1(\data_array.data1[13][12] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][12] ),
    .X(_04806_));
 sky130_fd_sc_hd__a221o_2 _07578_ (.A1(\data_array.data1[12][12] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][12] ),
    .C1(_04806_),
    .X(_04807_));
 sky130_fd_sc_hd__a22o_2 _07579_ (.A1(\data_array.data1[5][12] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][12] ),
    .X(_04808_));
 sky130_fd_sc_hd__a221o_2 _07580_ (.A1(\data_array.data1[4][12] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][12] ),
    .C1(_04808_),
    .X(_04809_));
 sky130_fd_sc_hd__a22o_2 _07581_ (.A1(_03506_),
    .A2(_04803_),
    .B1(_04807_),
    .B2(_03522_),
    .X(_04810_));
 sky130_fd_sc_hd__a22o_2 _07582_ (.A1(_03518_),
    .A2(_04805_),
    .B1(_04809_),
    .B2(_03526_),
    .X(_04811_));
 sky130_fd_sc_hd__or2_2 _07583_ (.A(_04810_),
    .B(_04811_),
    .X(_00067_));
 sky130_fd_sc_hd__a22o_2 _07584_ (.A1(\data_array.data1[13][13] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][13] ),
    .X(_04812_));
 sky130_fd_sc_hd__a221o_2 _07585_ (.A1(\data_array.data1[12][13] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][13] ),
    .C1(_04812_),
    .X(_04813_));
 sky130_fd_sc_hd__a22o_2 _07586_ (.A1(\data_array.data1[1][13] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][13] ),
    .X(_04814_));
 sky130_fd_sc_hd__a221o_2 _07587_ (.A1(\data_array.data1[0][13] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][13] ),
    .C1(_04814_),
    .X(_04815_));
 sky130_fd_sc_hd__a22o_2 _07588_ (.A1(\data_array.data1[9][13] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][13] ),
    .X(_04816_));
 sky130_fd_sc_hd__a221o_2 _07589_ (.A1(\data_array.data1[8][13] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][13] ),
    .C1(_04816_),
    .X(_04817_));
 sky130_fd_sc_hd__a22o_2 _07590_ (.A1(\data_array.data1[5][13] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][13] ),
    .X(_04818_));
 sky130_fd_sc_hd__a221o_2 _07591_ (.A1(\data_array.data1[4][13] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][13] ),
    .C1(_04818_),
    .X(_04819_));
 sky130_fd_sc_hd__a22o_2 _07592_ (.A1(_03522_),
    .A2(_04813_),
    .B1(_04817_),
    .B2(_03506_),
    .X(_04820_));
 sky130_fd_sc_hd__a22o_2 _07593_ (.A1(_03518_),
    .A2(_04815_),
    .B1(_04819_),
    .B2(_03526_),
    .X(_04821_));
 sky130_fd_sc_hd__or2_2 _07594_ (.A(_04820_),
    .B(_04821_),
    .X(_00068_));
 sky130_fd_sc_hd__a22o_2 _07595_ (.A1(\data_array.data1[9][14] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][14] ),
    .X(_04822_));
 sky130_fd_sc_hd__a221o_2 _07596_ (.A1(\data_array.data1[8][14] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][14] ),
    .C1(_04822_),
    .X(_04823_));
 sky130_fd_sc_hd__a22o_2 _07597_ (.A1(\data_array.data1[5][14] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][14] ),
    .X(_04824_));
 sky130_fd_sc_hd__a221o_2 _07598_ (.A1(\data_array.data1[4][14] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][14] ),
    .C1(_04824_),
    .X(_04825_));
 sky130_fd_sc_hd__a22o_2 _07599_ (.A1(\data_array.data1[13][14] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][14] ),
    .X(_04826_));
 sky130_fd_sc_hd__a221o_2 _07600_ (.A1(\data_array.data1[12][14] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][14] ),
    .C1(_04826_),
    .X(_04827_));
 sky130_fd_sc_hd__a22o_2 _07601_ (.A1(\data_array.data1[1][14] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][14] ),
    .X(_04828_));
 sky130_fd_sc_hd__a221o_2 _07602_ (.A1(\data_array.data1[0][14] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][14] ),
    .C1(_04828_),
    .X(_04829_));
 sky130_fd_sc_hd__a22o_2 _07603_ (.A1(_03506_),
    .A2(_04823_),
    .B1(_04827_),
    .B2(_03522_),
    .X(_04830_));
 sky130_fd_sc_hd__a22o_2 _07604_ (.A1(_03526_),
    .A2(_04825_),
    .B1(_04829_),
    .B2(_03518_),
    .X(_04831_));
 sky130_fd_sc_hd__or2_2 _07605_ (.A(_04830_),
    .B(_04831_),
    .X(_00069_));
 sky130_fd_sc_hd__a22o_2 _07606_ (.A1(\data_array.data1[9][15] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][15] ),
    .X(_04832_));
 sky130_fd_sc_hd__a221o_2 _07607_ (.A1(\data_array.data1[8][15] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][15] ),
    .C1(_04832_),
    .X(_04833_));
 sky130_fd_sc_hd__a22o_2 _07608_ (.A1(\data_array.data1[5][15] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][15] ),
    .X(_04834_));
 sky130_fd_sc_hd__a221o_2 _07609_ (.A1(\data_array.data1[4][15] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][15] ),
    .C1(_04834_),
    .X(_04835_));
 sky130_fd_sc_hd__a22o_2 _07610_ (.A1(\data_array.data1[13][15] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][15] ),
    .X(_04836_));
 sky130_fd_sc_hd__a221o_2 _07611_ (.A1(\data_array.data1[12][15] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][15] ),
    .C1(_04836_),
    .X(_04837_));
 sky130_fd_sc_hd__a22o_2 _07612_ (.A1(\data_array.data1[1][15] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][15] ),
    .X(_04838_));
 sky130_fd_sc_hd__a221o_2 _07613_ (.A1(\data_array.data1[0][15] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][15] ),
    .C1(_04838_),
    .X(_04839_));
 sky130_fd_sc_hd__a22o_2 _07614_ (.A1(_03506_),
    .A2(_04833_),
    .B1(_04837_),
    .B2(_03522_),
    .X(_04840_));
 sky130_fd_sc_hd__a22o_2 _07615_ (.A1(_03526_),
    .A2(_04835_),
    .B1(_04839_),
    .B2(_03518_),
    .X(_04841_));
 sky130_fd_sc_hd__or2_2 _07616_ (.A(_04840_),
    .B(_04841_),
    .X(_00070_));
 sky130_fd_sc_hd__a22o_2 _07617_ (.A1(\data_array.data1[9][16] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][16] ),
    .X(_04842_));
 sky130_fd_sc_hd__a221o_2 _07618_ (.A1(\data_array.data1[8][16] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][16] ),
    .C1(_04842_),
    .X(_04843_));
 sky130_fd_sc_hd__a22o_2 _07619_ (.A1(\data_array.data1[5][16] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][16] ),
    .X(_04844_));
 sky130_fd_sc_hd__a221o_2 _07620_ (.A1(\data_array.data1[4][16] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][16] ),
    .C1(_04844_),
    .X(_04845_));
 sky130_fd_sc_hd__a22o_2 _07621_ (.A1(\data_array.data1[13][16] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][16] ),
    .X(_04846_));
 sky130_fd_sc_hd__a221o_2 _07622_ (.A1(\data_array.data1[12][16] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][16] ),
    .C1(_04846_),
    .X(_04847_));
 sky130_fd_sc_hd__a22o_2 _07623_ (.A1(\data_array.data1[1][16] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][16] ),
    .X(_04848_));
 sky130_fd_sc_hd__a221o_2 _07624_ (.A1(\data_array.data1[0][16] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][16] ),
    .C1(_04848_),
    .X(_04849_));
 sky130_fd_sc_hd__a22o_2 _07625_ (.A1(_03506_),
    .A2(_04843_),
    .B1(_04847_),
    .B2(_03522_),
    .X(_04850_));
 sky130_fd_sc_hd__a22o_2 _07626_ (.A1(_03526_),
    .A2(_04845_),
    .B1(_04849_),
    .B2(_03518_),
    .X(_04851_));
 sky130_fd_sc_hd__or2_2 _07627_ (.A(_04850_),
    .B(_04851_),
    .X(_00071_));
 sky130_fd_sc_hd__a22o_2 _07628_ (.A1(\data_array.data1[13][17] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][17] ),
    .X(_04852_));
 sky130_fd_sc_hd__a221o_2 _07629_ (.A1(\data_array.data1[12][17] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][17] ),
    .C1(_04852_),
    .X(_04853_));
 sky130_fd_sc_hd__a22o_2 _07630_ (.A1(\data_array.data1[1][17] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][17] ),
    .X(_04854_));
 sky130_fd_sc_hd__a221o_2 _07631_ (.A1(\data_array.data1[0][17] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][17] ),
    .C1(_04854_),
    .X(_04855_));
 sky130_fd_sc_hd__a22o_2 _07632_ (.A1(\data_array.data1[9][17] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][17] ),
    .X(_04856_));
 sky130_fd_sc_hd__a221o_2 _07633_ (.A1(\data_array.data1[8][17] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][17] ),
    .C1(_04856_),
    .X(_04857_));
 sky130_fd_sc_hd__a22o_2 _07634_ (.A1(\data_array.data1[5][17] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][17] ),
    .X(_04858_));
 sky130_fd_sc_hd__a221o_2 _07635_ (.A1(\data_array.data1[4][17] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][17] ),
    .C1(_04858_),
    .X(_04859_));
 sky130_fd_sc_hd__a22o_2 _07636_ (.A1(_03522_),
    .A2(_04853_),
    .B1(_04857_),
    .B2(_03506_),
    .X(_04860_));
 sky130_fd_sc_hd__a22o_2 _07637_ (.A1(_03518_),
    .A2(_04855_),
    .B1(_04859_),
    .B2(_03526_),
    .X(_04861_));
 sky130_fd_sc_hd__or2_2 _07638_ (.A(_04860_),
    .B(_04861_),
    .X(_00072_));
 sky130_fd_sc_hd__a22o_2 _07639_ (.A1(\data_array.data1[9][18] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][18] ),
    .X(_04862_));
 sky130_fd_sc_hd__a221o_2 _07640_ (.A1(\data_array.data1[8][18] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][18] ),
    .C1(_04862_),
    .X(_04863_));
 sky130_fd_sc_hd__a22o_2 _07641_ (.A1(\data_array.data1[5][18] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][18] ),
    .X(_04864_));
 sky130_fd_sc_hd__a221o_2 _07642_ (.A1(\data_array.data1[4][18] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][18] ),
    .C1(_04864_),
    .X(_04865_));
 sky130_fd_sc_hd__a22o_2 _07643_ (.A1(\data_array.data1[13][18] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][18] ),
    .X(_04866_));
 sky130_fd_sc_hd__a221o_2 _07644_ (.A1(\data_array.data1[12][18] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][18] ),
    .C1(_04866_),
    .X(_04867_));
 sky130_fd_sc_hd__a22o_2 _07645_ (.A1(\data_array.data1[1][18] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][18] ),
    .X(_04868_));
 sky130_fd_sc_hd__a221o_2 _07646_ (.A1(\data_array.data1[0][18] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][18] ),
    .C1(_04868_),
    .X(_04869_));
 sky130_fd_sc_hd__a22o_2 _07647_ (.A1(_03506_),
    .A2(_04863_),
    .B1(_04867_),
    .B2(_03522_),
    .X(_04870_));
 sky130_fd_sc_hd__a22o_2 _07648_ (.A1(_03526_),
    .A2(_04865_),
    .B1(_04869_),
    .B2(_03518_),
    .X(_04871_));
 sky130_fd_sc_hd__or2_2 _07649_ (.A(_04870_),
    .B(_04871_),
    .X(_00073_));
 sky130_fd_sc_hd__a22o_2 _07650_ (.A1(\data_array.data1[13][19] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][19] ),
    .X(_04872_));
 sky130_fd_sc_hd__a221o_2 _07651_ (.A1(\data_array.data1[12][19] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][19] ),
    .C1(_04872_),
    .X(_04873_));
 sky130_fd_sc_hd__a22o_2 _07652_ (.A1(\data_array.data1[5][19] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][19] ),
    .X(_04874_));
 sky130_fd_sc_hd__a221o_2 _07653_ (.A1(\data_array.data1[4][19] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][19] ),
    .C1(_04874_),
    .X(_04875_));
 sky130_fd_sc_hd__a22o_2 _07654_ (.A1(\data_array.data1[9][19] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][19] ),
    .X(_04876_));
 sky130_fd_sc_hd__a221o_2 _07655_ (.A1(\data_array.data1[8][19] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][19] ),
    .C1(_04876_),
    .X(_04877_));
 sky130_fd_sc_hd__a22o_2 _07656_ (.A1(\data_array.data1[1][19] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][19] ),
    .X(_04878_));
 sky130_fd_sc_hd__a221o_2 _07657_ (.A1(\data_array.data1[0][19] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][19] ),
    .C1(_04878_),
    .X(_04879_));
 sky130_fd_sc_hd__a22o_2 _07658_ (.A1(_03522_),
    .A2(_04873_),
    .B1(_04877_),
    .B2(_03506_),
    .X(_04880_));
 sky130_fd_sc_hd__a22o_2 _07659_ (.A1(_03526_),
    .A2(_04875_),
    .B1(_04879_),
    .B2(_03518_),
    .X(_04881_));
 sky130_fd_sc_hd__or2_2 _07660_ (.A(_04880_),
    .B(_04881_),
    .X(_00074_));
 sky130_fd_sc_hd__a22o_2 _07661_ (.A1(\data_array.data1[13][20] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][20] ),
    .X(_04882_));
 sky130_fd_sc_hd__a221o_2 _07662_ (.A1(\data_array.data1[12][20] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][20] ),
    .C1(_04882_),
    .X(_04883_));
 sky130_fd_sc_hd__a22o_2 _07663_ (.A1(\data_array.data1[5][20] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][20] ),
    .X(_04884_));
 sky130_fd_sc_hd__a221o_2 _07664_ (.A1(\data_array.data1[4][20] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][20] ),
    .C1(_04884_),
    .X(_04885_));
 sky130_fd_sc_hd__a22o_2 _07665_ (.A1(\data_array.data1[9][20] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][20] ),
    .X(_04886_));
 sky130_fd_sc_hd__a221o_2 _07666_ (.A1(\data_array.data1[8][20] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][20] ),
    .C1(_04886_),
    .X(_04887_));
 sky130_fd_sc_hd__a22o_2 _07667_ (.A1(\data_array.data1[1][20] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][20] ),
    .X(_04888_));
 sky130_fd_sc_hd__a221o_2 _07668_ (.A1(\data_array.data1[0][20] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][20] ),
    .C1(_04888_),
    .X(_04889_));
 sky130_fd_sc_hd__a22o_2 _07669_ (.A1(_03522_),
    .A2(_04883_),
    .B1(_04887_),
    .B2(_03506_),
    .X(_04890_));
 sky130_fd_sc_hd__a22o_2 _07670_ (.A1(_03526_),
    .A2(_04885_),
    .B1(_04889_),
    .B2(_03518_),
    .X(_04891_));
 sky130_fd_sc_hd__or2_2 _07671_ (.A(_04890_),
    .B(_04891_),
    .X(_00076_));
 sky130_fd_sc_hd__a22o_2 _07672_ (.A1(\data_array.data1[9][21] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][21] ),
    .X(_04892_));
 sky130_fd_sc_hd__a221o_2 _07673_ (.A1(\data_array.data1[8][21] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][21] ),
    .C1(_04892_),
    .X(_04893_));
 sky130_fd_sc_hd__a22o_2 _07674_ (.A1(\data_array.data1[1][21] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][21] ),
    .X(_04894_));
 sky130_fd_sc_hd__a221o_2 _07675_ (.A1(\data_array.data1[0][21] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][21] ),
    .C1(_04894_),
    .X(_04895_));
 sky130_fd_sc_hd__a22o_2 _07676_ (.A1(\data_array.data1[13][21] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][21] ),
    .X(_04896_));
 sky130_fd_sc_hd__a221o_2 _07677_ (.A1(\data_array.data1[12][21] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][21] ),
    .C1(_04896_),
    .X(_04897_));
 sky130_fd_sc_hd__a22o_2 _07678_ (.A1(\data_array.data1[5][21] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][21] ),
    .X(_04898_));
 sky130_fd_sc_hd__a221o_2 _07679_ (.A1(\data_array.data1[4][21] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][21] ),
    .C1(_04898_),
    .X(_04899_));
 sky130_fd_sc_hd__a22o_2 _07680_ (.A1(_03506_),
    .A2(_04893_),
    .B1(_04897_),
    .B2(_03522_),
    .X(_04900_));
 sky130_fd_sc_hd__a22o_2 _07681_ (.A1(_03518_),
    .A2(_04895_),
    .B1(_04899_),
    .B2(_03526_),
    .X(_04901_));
 sky130_fd_sc_hd__or2_2 _07682_ (.A(_04900_),
    .B(_04901_),
    .X(_00077_));
 sky130_fd_sc_hd__a22o_2 _07683_ (.A1(\data_array.data1[9][22] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][22] ),
    .X(_04902_));
 sky130_fd_sc_hd__a221o_2 _07684_ (.A1(\data_array.data1[8][22] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][22] ),
    .C1(_04902_),
    .X(_04903_));
 sky130_fd_sc_hd__a22o_2 _07685_ (.A1(\data_array.data1[1][22] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][22] ),
    .X(_04904_));
 sky130_fd_sc_hd__a221o_2 _07686_ (.A1(\data_array.data1[0][22] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][22] ),
    .C1(_04904_),
    .X(_04905_));
 sky130_fd_sc_hd__a22o_2 _07687_ (.A1(\data_array.data1[13][22] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][22] ),
    .X(_04906_));
 sky130_fd_sc_hd__a221o_2 _07688_ (.A1(\data_array.data1[12][22] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][22] ),
    .C1(_04906_),
    .X(_04907_));
 sky130_fd_sc_hd__a22o_2 _07689_ (.A1(\data_array.data1[5][22] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][22] ),
    .X(_04908_));
 sky130_fd_sc_hd__a221o_2 _07690_ (.A1(\data_array.data1[4][22] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][22] ),
    .C1(_04908_),
    .X(_04909_));
 sky130_fd_sc_hd__a22o_2 _07691_ (.A1(_03506_),
    .A2(_04903_),
    .B1(_04907_),
    .B2(_03522_),
    .X(_04910_));
 sky130_fd_sc_hd__a22o_2 _07692_ (.A1(_03518_),
    .A2(_04905_),
    .B1(_04909_),
    .B2(_03526_),
    .X(_04911_));
 sky130_fd_sc_hd__or2_2 _07693_ (.A(_04910_),
    .B(_04911_),
    .X(_00078_));
 sky130_fd_sc_hd__a22o_2 _07694_ (.A1(\data_array.data1[13][23] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][23] ),
    .X(_04912_));
 sky130_fd_sc_hd__a221o_2 _07695_ (.A1(\data_array.data1[12][23] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][23] ),
    .C1(_04912_),
    .X(_04913_));
 sky130_fd_sc_hd__a22o_2 _07696_ (.A1(\data_array.data1[1][23] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][23] ),
    .X(_04914_));
 sky130_fd_sc_hd__a221o_2 _07697_ (.A1(\data_array.data1[0][23] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][23] ),
    .C1(_04914_),
    .X(_04915_));
 sky130_fd_sc_hd__a22o_2 _07698_ (.A1(\data_array.data1[9][23] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][23] ),
    .X(_04916_));
 sky130_fd_sc_hd__a221o_2 _07699_ (.A1(\data_array.data1[8][23] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][23] ),
    .C1(_04916_),
    .X(_04917_));
 sky130_fd_sc_hd__a22o_2 _07700_ (.A1(\data_array.data1[5][23] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][23] ),
    .X(_04918_));
 sky130_fd_sc_hd__a221o_2 _07701_ (.A1(\data_array.data1[4][23] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][23] ),
    .C1(_04918_),
    .X(_04919_));
 sky130_fd_sc_hd__a22o_2 _07702_ (.A1(_03522_),
    .A2(_04913_),
    .B1(_04917_),
    .B2(_03506_),
    .X(_04920_));
 sky130_fd_sc_hd__a22o_2 _07703_ (.A1(_03518_),
    .A2(_04915_),
    .B1(_04919_),
    .B2(_03526_),
    .X(_04921_));
 sky130_fd_sc_hd__or2_2 _07704_ (.A(_04920_),
    .B(_04921_),
    .X(_00079_));
 sky130_fd_sc_hd__a22o_2 _07705_ (.A1(\data_array.data1[13][24] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][24] ),
    .X(_04922_));
 sky130_fd_sc_hd__a221o_2 _07706_ (.A1(\data_array.data1[12][24] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][24] ),
    .C1(_04922_),
    .X(_04923_));
 sky130_fd_sc_hd__a22o_2 _07707_ (.A1(\data_array.data1[5][24] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][24] ),
    .X(_04924_));
 sky130_fd_sc_hd__a221o_2 _07708_ (.A1(\data_array.data1[4][24] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][24] ),
    .C1(_04924_),
    .X(_04925_));
 sky130_fd_sc_hd__a22o_2 _07709_ (.A1(\data_array.data1[9][24] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][24] ),
    .X(_04926_));
 sky130_fd_sc_hd__a221o_2 _07710_ (.A1(\data_array.data1[8][24] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][24] ),
    .C1(_04926_),
    .X(_04927_));
 sky130_fd_sc_hd__a22o_2 _07711_ (.A1(\data_array.data1[1][24] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][24] ),
    .X(_04928_));
 sky130_fd_sc_hd__a221o_2 _07712_ (.A1(\data_array.data1[0][24] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][24] ),
    .C1(_04928_),
    .X(_04929_));
 sky130_fd_sc_hd__a22o_2 _07713_ (.A1(_03522_),
    .A2(_04923_),
    .B1(_04927_),
    .B2(_03506_),
    .X(_04930_));
 sky130_fd_sc_hd__a22o_2 _07714_ (.A1(_03526_),
    .A2(_04925_),
    .B1(_04929_),
    .B2(_03518_),
    .X(_04931_));
 sky130_fd_sc_hd__or2_2 _07715_ (.A(_04930_),
    .B(_04931_),
    .X(_00080_));
 sky130_fd_sc_hd__a22o_2 _07716_ (.A1(\data_array.data1[13][25] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][25] ),
    .X(_04932_));
 sky130_fd_sc_hd__a221o_2 _07717_ (.A1(\data_array.data1[12][25] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][25] ),
    .C1(_04932_),
    .X(_04933_));
 sky130_fd_sc_hd__a22o_2 _07718_ (.A1(\data_array.data1[1][25] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][25] ),
    .X(_04934_));
 sky130_fd_sc_hd__a221o_2 _07719_ (.A1(\data_array.data1[0][25] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][25] ),
    .C1(_04934_),
    .X(_04935_));
 sky130_fd_sc_hd__a22o_2 _07720_ (.A1(\data_array.data1[9][25] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][25] ),
    .X(_04936_));
 sky130_fd_sc_hd__a221o_2 _07721_ (.A1(\data_array.data1[8][25] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][25] ),
    .C1(_04936_),
    .X(_04937_));
 sky130_fd_sc_hd__a22o_2 _07722_ (.A1(\data_array.data1[5][25] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][25] ),
    .X(_04938_));
 sky130_fd_sc_hd__a221o_2 _07723_ (.A1(\data_array.data1[4][25] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][25] ),
    .C1(_04938_),
    .X(_04939_));
 sky130_fd_sc_hd__a22o_2 _07724_ (.A1(_03522_),
    .A2(_04933_),
    .B1(_04937_),
    .B2(_03506_),
    .X(_04940_));
 sky130_fd_sc_hd__a22o_2 _07725_ (.A1(_03518_),
    .A2(_04935_),
    .B1(_04939_),
    .B2(_03526_),
    .X(_04941_));
 sky130_fd_sc_hd__or2_2 _07726_ (.A(_04940_),
    .B(_04941_),
    .X(_00081_));
 sky130_fd_sc_hd__a22o_2 _07727_ (.A1(\data_array.data1[9][26] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][26] ),
    .X(_04942_));
 sky130_fd_sc_hd__a221o_2 _07728_ (.A1(\data_array.data1[8][26] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][26] ),
    .C1(_04942_),
    .X(_04943_));
 sky130_fd_sc_hd__a22o_2 _07729_ (.A1(\data_array.data1[5][26] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][26] ),
    .X(_04944_));
 sky130_fd_sc_hd__a221o_2 _07730_ (.A1(\data_array.data1[4][26] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][26] ),
    .C1(_04944_),
    .X(_04945_));
 sky130_fd_sc_hd__a22o_2 _07731_ (.A1(\data_array.data1[13][26] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][26] ),
    .X(_04946_));
 sky130_fd_sc_hd__a221o_2 _07732_ (.A1(\data_array.data1[12][26] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][26] ),
    .C1(_04946_),
    .X(_04947_));
 sky130_fd_sc_hd__a22o_2 _07733_ (.A1(\data_array.data1[1][26] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][26] ),
    .X(_04948_));
 sky130_fd_sc_hd__a221o_2 _07734_ (.A1(\data_array.data1[0][26] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][26] ),
    .C1(_04948_),
    .X(_04949_));
 sky130_fd_sc_hd__a22o_2 _07735_ (.A1(_03506_),
    .A2(_04943_),
    .B1(_04947_),
    .B2(_03522_),
    .X(_04950_));
 sky130_fd_sc_hd__a22o_2 _07736_ (.A1(_03526_),
    .A2(_04945_),
    .B1(_04949_),
    .B2(_03518_),
    .X(_04951_));
 sky130_fd_sc_hd__or2_2 _07737_ (.A(_04950_),
    .B(_04951_),
    .X(_00082_));
 sky130_fd_sc_hd__a22o_2 _07738_ (.A1(\data_array.data1[9][27] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][27] ),
    .X(_04952_));
 sky130_fd_sc_hd__a221o_2 _07739_ (.A1(\data_array.data1[8][27] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][27] ),
    .C1(_04952_),
    .X(_04953_));
 sky130_fd_sc_hd__a22o_2 _07740_ (.A1(\data_array.data1[1][27] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][27] ),
    .X(_04954_));
 sky130_fd_sc_hd__a221o_2 _07741_ (.A1(\data_array.data1[0][27] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][27] ),
    .C1(_04954_),
    .X(_04955_));
 sky130_fd_sc_hd__a22o_2 _07742_ (.A1(\data_array.data1[13][27] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][27] ),
    .X(_04956_));
 sky130_fd_sc_hd__a221o_2 _07743_ (.A1(\data_array.data1[12][27] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][27] ),
    .C1(_04956_),
    .X(_04957_));
 sky130_fd_sc_hd__a22o_2 _07744_ (.A1(\data_array.data1[5][27] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][27] ),
    .X(_04958_));
 sky130_fd_sc_hd__a221o_2 _07745_ (.A1(\data_array.data1[4][27] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][27] ),
    .C1(_04958_),
    .X(_04959_));
 sky130_fd_sc_hd__a22o_2 _07746_ (.A1(_03506_),
    .A2(_04953_),
    .B1(_04957_),
    .B2(_03522_),
    .X(_04960_));
 sky130_fd_sc_hd__a22o_2 _07747_ (.A1(_03518_),
    .A2(_04955_),
    .B1(_04959_),
    .B2(_03526_),
    .X(_04961_));
 sky130_fd_sc_hd__or2_2 _07748_ (.A(_04960_),
    .B(_04961_),
    .X(_00083_));
 sky130_fd_sc_hd__a22o_2 _07749_ (.A1(\data_array.data1[9][28] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][28] ),
    .X(_04962_));
 sky130_fd_sc_hd__a221o_2 _07750_ (.A1(\data_array.data1[8][28] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][28] ),
    .C1(_04962_),
    .X(_04963_));
 sky130_fd_sc_hd__a22o_2 _07751_ (.A1(\data_array.data1[5][28] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][28] ),
    .X(_04964_));
 sky130_fd_sc_hd__a221o_2 _07752_ (.A1(\data_array.data1[4][28] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][28] ),
    .C1(_04964_),
    .X(_04965_));
 sky130_fd_sc_hd__a22o_2 _07753_ (.A1(\data_array.data1[13][28] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][28] ),
    .X(_04966_));
 sky130_fd_sc_hd__a221o_2 _07754_ (.A1(\data_array.data1[12][28] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][28] ),
    .C1(_04966_),
    .X(_04967_));
 sky130_fd_sc_hd__a22o_2 _07755_ (.A1(\data_array.data1[1][28] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][28] ),
    .X(_04968_));
 sky130_fd_sc_hd__a221o_2 _07756_ (.A1(\data_array.data1[0][28] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][28] ),
    .C1(_04968_),
    .X(_04969_));
 sky130_fd_sc_hd__a22o_2 _07757_ (.A1(_03506_),
    .A2(_04963_),
    .B1(_04967_),
    .B2(_03522_),
    .X(_04970_));
 sky130_fd_sc_hd__a22o_2 _07758_ (.A1(_03526_),
    .A2(_04965_),
    .B1(_04969_),
    .B2(_03518_),
    .X(_04971_));
 sky130_fd_sc_hd__or2_2 _07759_ (.A(_04970_),
    .B(_04971_),
    .X(_00084_));
 sky130_fd_sc_hd__a22o_2 _07760_ (.A1(\data_array.data1[13][29] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][29] ),
    .X(_04972_));
 sky130_fd_sc_hd__a221o_2 _07761_ (.A1(\data_array.data1[12][29] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][29] ),
    .C1(_04972_),
    .X(_04973_));
 sky130_fd_sc_hd__a22o_2 _07762_ (.A1(\data_array.data1[1][29] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][29] ),
    .X(_04974_));
 sky130_fd_sc_hd__a221o_2 _07763_ (.A1(\data_array.data1[0][29] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][29] ),
    .C1(_04974_),
    .X(_04975_));
 sky130_fd_sc_hd__a22o_2 _07764_ (.A1(\data_array.data1[9][29] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][29] ),
    .X(_04976_));
 sky130_fd_sc_hd__a221o_2 _07765_ (.A1(\data_array.data1[8][29] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][29] ),
    .C1(_04976_),
    .X(_04977_));
 sky130_fd_sc_hd__a22o_2 _07766_ (.A1(\data_array.data1[5][29] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][29] ),
    .X(_04978_));
 sky130_fd_sc_hd__a221o_2 _07767_ (.A1(\data_array.data1[4][29] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][29] ),
    .C1(_04978_),
    .X(_04979_));
 sky130_fd_sc_hd__a22o_2 _07768_ (.A1(_03522_),
    .A2(_04973_),
    .B1(_04977_),
    .B2(_03506_),
    .X(_04980_));
 sky130_fd_sc_hd__a22o_2 _07769_ (.A1(_03518_),
    .A2(_04975_),
    .B1(_04979_),
    .B2(_03526_),
    .X(_04981_));
 sky130_fd_sc_hd__or2_2 _07770_ (.A(_04980_),
    .B(_04981_),
    .X(_00085_));
 sky130_fd_sc_hd__a22o_2 _07771_ (.A1(\data_array.data1[9][30] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][30] ),
    .X(_04982_));
 sky130_fd_sc_hd__a221o_2 _07772_ (.A1(\data_array.data1[8][30] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][30] ),
    .C1(_04982_),
    .X(_04983_));
 sky130_fd_sc_hd__a22o_2 _07773_ (.A1(\data_array.data1[5][30] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][30] ),
    .X(_04984_));
 sky130_fd_sc_hd__a221o_2 _07774_ (.A1(\data_array.data1[4][30] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][30] ),
    .C1(_04984_),
    .X(_04985_));
 sky130_fd_sc_hd__a22o_2 _07775_ (.A1(\data_array.data1[13][30] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][30] ),
    .X(_04986_));
 sky130_fd_sc_hd__a221o_2 _07776_ (.A1(\data_array.data1[12][30] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][30] ),
    .C1(_04986_),
    .X(_04987_));
 sky130_fd_sc_hd__a22o_2 _07777_ (.A1(\data_array.data1[1][30] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][30] ),
    .X(_04988_));
 sky130_fd_sc_hd__a221o_2 _07778_ (.A1(\data_array.data1[0][30] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][30] ),
    .C1(_04988_),
    .X(_04989_));
 sky130_fd_sc_hd__a22o_2 _07779_ (.A1(_03506_),
    .A2(_04983_),
    .B1(_04987_),
    .B2(_03522_),
    .X(_04990_));
 sky130_fd_sc_hd__a22o_2 _07780_ (.A1(_03526_),
    .A2(_04985_),
    .B1(_04989_),
    .B2(_03518_),
    .X(_04991_));
 sky130_fd_sc_hd__or2_2 _07781_ (.A(_04990_),
    .B(_04991_),
    .X(_00087_));
 sky130_fd_sc_hd__a22o_2 _07782_ (.A1(\data_array.data1[13][31] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][31] ),
    .X(_04992_));
 sky130_fd_sc_hd__a221o_2 _07783_ (.A1(\data_array.data1[12][31] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][31] ),
    .C1(_04992_),
    .X(_04993_));
 sky130_fd_sc_hd__a22o_2 _07784_ (.A1(\data_array.data1[5][31] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][31] ),
    .X(_04994_));
 sky130_fd_sc_hd__a221o_2 _07785_ (.A1(\data_array.data1[4][31] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][31] ),
    .C1(_04994_),
    .X(_04995_));
 sky130_fd_sc_hd__a22o_2 _07786_ (.A1(\data_array.data1[9][31] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][31] ),
    .X(_04996_));
 sky130_fd_sc_hd__a221o_2 _07787_ (.A1(\data_array.data1[8][31] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][31] ),
    .C1(_04996_),
    .X(_04997_));
 sky130_fd_sc_hd__a22o_2 _07788_ (.A1(\data_array.data1[1][31] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][31] ),
    .X(_04998_));
 sky130_fd_sc_hd__a221o_2 _07789_ (.A1(\data_array.data1[0][31] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][31] ),
    .C1(_04998_),
    .X(_04999_));
 sky130_fd_sc_hd__a22o_2 _07790_ (.A1(_03522_),
    .A2(_04993_),
    .B1(_04997_),
    .B2(_03506_),
    .X(_05000_));
 sky130_fd_sc_hd__a22o_2 _07791_ (.A1(_03526_),
    .A2(_04995_),
    .B1(_04999_),
    .B2(_03518_),
    .X(_05001_));
 sky130_fd_sc_hd__or2_2 _07792_ (.A(_05000_),
    .B(_05001_),
    .X(_00088_));
 sky130_fd_sc_hd__a22o_2 _07793_ (.A1(\data_array.data1[13][32] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][32] ),
    .X(_05002_));
 sky130_fd_sc_hd__a221o_2 _07794_ (.A1(\data_array.data1[12][32] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][32] ),
    .C1(_05002_),
    .X(_05003_));
 sky130_fd_sc_hd__a22o_2 _07795_ (.A1(\data_array.data1[1][32] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][32] ),
    .X(_05004_));
 sky130_fd_sc_hd__a221o_2 _07796_ (.A1(\data_array.data1[0][32] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][32] ),
    .C1(_05004_),
    .X(_05005_));
 sky130_fd_sc_hd__a22o_2 _07797_ (.A1(\data_array.data1[9][32] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][32] ),
    .X(_05006_));
 sky130_fd_sc_hd__a221o_2 _07798_ (.A1(\data_array.data1[8][32] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][32] ),
    .C1(_05006_),
    .X(_05007_));
 sky130_fd_sc_hd__a22o_2 _07799_ (.A1(\data_array.data1[5][32] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][32] ),
    .X(_05008_));
 sky130_fd_sc_hd__a221o_2 _07800_ (.A1(\data_array.data1[4][32] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][32] ),
    .C1(_05008_),
    .X(_05009_));
 sky130_fd_sc_hd__a22o_2 _07801_ (.A1(_03522_),
    .A2(_05003_),
    .B1(_05007_),
    .B2(_03506_),
    .X(_05010_));
 sky130_fd_sc_hd__a22o_2 _07802_ (.A1(_03518_),
    .A2(_05005_),
    .B1(_05009_),
    .B2(_03526_),
    .X(_05011_));
 sky130_fd_sc_hd__or2_2 _07803_ (.A(_05010_),
    .B(_05011_),
    .X(_00089_));
 sky130_fd_sc_hd__a22o_2 _07804_ (.A1(\data_array.data1[13][33] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][33] ),
    .X(_05012_));
 sky130_fd_sc_hd__a221o_2 _07805_ (.A1(\data_array.data1[12][33] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][33] ),
    .C1(_05012_),
    .X(_05013_));
 sky130_fd_sc_hd__a22o_2 _07806_ (.A1(\data_array.data1[1][33] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][33] ),
    .X(_05014_));
 sky130_fd_sc_hd__a221o_2 _07807_ (.A1(\data_array.data1[0][33] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][33] ),
    .C1(_05014_),
    .X(_05015_));
 sky130_fd_sc_hd__a22o_2 _07808_ (.A1(\data_array.data1[9][33] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][33] ),
    .X(_05016_));
 sky130_fd_sc_hd__a221o_2 _07809_ (.A1(\data_array.data1[8][33] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][33] ),
    .C1(_05016_),
    .X(_05017_));
 sky130_fd_sc_hd__a22o_2 _07810_ (.A1(\data_array.data1[5][33] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][33] ),
    .X(_05018_));
 sky130_fd_sc_hd__a221o_2 _07811_ (.A1(\data_array.data1[4][33] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][33] ),
    .C1(_05018_),
    .X(_05019_));
 sky130_fd_sc_hd__a22o_2 _07812_ (.A1(_03522_),
    .A2(_05013_),
    .B1(_05017_),
    .B2(_03506_),
    .X(_05020_));
 sky130_fd_sc_hd__a22o_2 _07813_ (.A1(_03518_),
    .A2(_05015_),
    .B1(_05019_),
    .B2(_03526_),
    .X(_05021_));
 sky130_fd_sc_hd__or2_2 _07814_ (.A(_05020_),
    .B(_05021_),
    .X(_00090_));
 sky130_fd_sc_hd__a22o_2 _07815_ (.A1(\data_array.data1[13][34] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][34] ),
    .X(_05022_));
 sky130_fd_sc_hd__a221o_2 _07816_ (.A1(\data_array.data1[12][34] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][34] ),
    .C1(_05022_),
    .X(_05023_));
 sky130_fd_sc_hd__a22o_2 _07817_ (.A1(\data_array.data1[5][34] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][34] ),
    .X(_05024_));
 sky130_fd_sc_hd__a221o_2 _07818_ (.A1(\data_array.data1[4][34] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][34] ),
    .C1(_05024_),
    .X(_05025_));
 sky130_fd_sc_hd__a22o_2 _07819_ (.A1(\data_array.data1[9][34] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][34] ),
    .X(_05026_));
 sky130_fd_sc_hd__a221o_2 _07820_ (.A1(\data_array.data1[8][34] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][34] ),
    .C1(_05026_),
    .X(_05027_));
 sky130_fd_sc_hd__a22o_2 _07821_ (.A1(\data_array.data1[1][34] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][34] ),
    .X(_05028_));
 sky130_fd_sc_hd__a221o_2 _07822_ (.A1(\data_array.data1[0][34] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][34] ),
    .C1(_05028_),
    .X(_05029_));
 sky130_fd_sc_hd__a22o_2 _07823_ (.A1(_03522_),
    .A2(_05023_),
    .B1(_05027_),
    .B2(_03506_),
    .X(_05030_));
 sky130_fd_sc_hd__a22o_2 _07824_ (.A1(_03526_),
    .A2(_05025_),
    .B1(_05029_),
    .B2(_03518_),
    .X(_05031_));
 sky130_fd_sc_hd__or2_2 _07825_ (.A(_05030_),
    .B(_05031_),
    .X(_00091_));
 sky130_fd_sc_hd__a22o_2 _07826_ (.A1(\data_array.data1[13][35] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][35] ),
    .X(_05032_));
 sky130_fd_sc_hd__a221o_2 _07827_ (.A1(\data_array.data1[12][35] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][35] ),
    .C1(_05032_),
    .X(_05033_));
 sky130_fd_sc_hd__a22o_2 _07828_ (.A1(\data_array.data1[5][35] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][35] ),
    .X(_05034_));
 sky130_fd_sc_hd__a221o_2 _07829_ (.A1(\data_array.data1[4][35] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][35] ),
    .C1(_05034_),
    .X(_05035_));
 sky130_fd_sc_hd__a22o_2 _07830_ (.A1(\data_array.data1[9][35] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][35] ),
    .X(_05036_));
 sky130_fd_sc_hd__a221o_2 _07831_ (.A1(\data_array.data1[8][35] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][35] ),
    .C1(_05036_),
    .X(_05037_));
 sky130_fd_sc_hd__a22o_2 _07832_ (.A1(\data_array.data1[1][35] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][35] ),
    .X(_05038_));
 sky130_fd_sc_hd__a221o_2 _07833_ (.A1(\data_array.data1[0][35] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][35] ),
    .C1(_05038_),
    .X(_05039_));
 sky130_fd_sc_hd__a22o_2 _07834_ (.A1(_03522_),
    .A2(_05033_),
    .B1(_05037_),
    .B2(_03506_),
    .X(_05040_));
 sky130_fd_sc_hd__a22o_2 _07835_ (.A1(_03526_),
    .A2(_05035_),
    .B1(_05039_),
    .B2(_03518_),
    .X(_05041_));
 sky130_fd_sc_hd__or2_2 _07836_ (.A(_05040_),
    .B(_05041_),
    .X(_00092_));
 sky130_fd_sc_hd__a22o_2 _07837_ (.A1(\data_array.data1[9][36] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][36] ),
    .X(_05042_));
 sky130_fd_sc_hd__a221o_2 _07838_ (.A1(\data_array.data1[8][36] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][36] ),
    .C1(_05042_),
    .X(_05043_));
 sky130_fd_sc_hd__a22o_2 _07839_ (.A1(\data_array.data1[5][36] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][36] ),
    .X(_05044_));
 sky130_fd_sc_hd__a221o_2 _07840_ (.A1(\data_array.data1[4][36] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][36] ),
    .C1(_05044_),
    .X(_05045_));
 sky130_fd_sc_hd__a22o_2 _07841_ (.A1(\data_array.data1[13][36] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][36] ),
    .X(_05046_));
 sky130_fd_sc_hd__a221o_2 _07842_ (.A1(\data_array.data1[12][36] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][36] ),
    .C1(_05046_),
    .X(_05047_));
 sky130_fd_sc_hd__a22o_2 _07843_ (.A1(\data_array.data1[1][36] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][36] ),
    .X(_05048_));
 sky130_fd_sc_hd__a221o_2 _07844_ (.A1(\data_array.data1[0][36] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][36] ),
    .C1(_05048_),
    .X(_05049_));
 sky130_fd_sc_hd__a22o_2 _07845_ (.A1(_03506_),
    .A2(_05043_),
    .B1(_05047_),
    .B2(_03522_),
    .X(_05050_));
 sky130_fd_sc_hd__a22o_2 _07846_ (.A1(_03526_),
    .A2(_05045_),
    .B1(_05049_),
    .B2(_03518_),
    .X(_05051_));
 sky130_fd_sc_hd__or2_2 _07847_ (.A(_05050_),
    .B(_05051_),
    .X(_00093_));
 sky130_fd_sc_hd__a22o_2 _07848_ (.A1(\data_array.data1[9][37] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][37] ),
    .X(_05052_));
 sky130_fd_sc_hd__a221o_2 _07849_ (.A1(\data_array.data1[8][37] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][37] ),
    .C1(_05052_),
    .X(_05053_));
 sky130_fd_sc_hd__a22o_2 _07850_ (.A1(\data_array.data1[1][37] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][37] ),
    .X(_05054_));
 sky130_fd_sc_hd__a221o_2 _07851_ (.A1(\data_array.data1[0][37] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][37] ),
    .C1(_05054_),
    .X(_05055_));
 sky130_fd_sc_hd__a22o_2 _07852_ (.A1(\data_array.data1[13][37] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][37] ),
    .X(_05056_));
 sky130_fd_sc_hd__a221o_2 _07853_ (.A1(\data_array.data1[12][37] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][37] ),
    .C1(_05056_),
    .X(_05057_));
 sky130_fd_sc_hd__a22o_2 _07854_ (.A1(\data_array.data1[5][37] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][37] ),
    .X(_05058_));
 sky130_fd_sc_hd__a221o_2 _07855_ (.A1(\data_array.data1[4][37] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][37] ),
    .C1(_05058_),
    .X(_05059_));
 sky130_fd_sc_hd__a22o_2 _07856_ (.A1(_03506_),
    .A2(_05053_),
    .B1(_05057_),
    .B2(_03522_),
    .X(_05060_));
 sky130_fd_sc_hd__a22o_2 _07857_ (.A1(_03518_),
    .A2(_05055_),
    .B1(_05059_),
    .B2(_03526_),
    .X(_05061_));
 sky130_fd_sc_hd__or2_2 _07858_ (.A(_05060_),
    .B(_05061_),
    .X(_00094_));
 sky130_fd_sc_hd__a22o_2 _07859_ (.A1(\data_array.data1[9][38] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][38] ),
    .X(_05062_));
 sky130_fd_sc_hd__a221o_2 _07860_ (.A1(\data_array.data1[8][38] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][38] ),
    .C1(_05062_),
    .X(_05063_));
 sky130_fd_sc_hd__a22o_2 _07861_ (.A1(\data_array.data1[1][38] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][38] ),
    .X(_05064_));
 sky130_fd_sc_hd__a221o_2 _07862_ (.A1(\data_array.data1[0][38] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][38] ),
    .C1(_05064_),
    .X(_05065_));
 sky130_fd_sc_hd__a22o_2 _07863_ (.A1(\data_array.data1[13][38] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][38] ),
    .X(_05066_));
 sky130_fd_sc_hd__a221o_2 _07864_ (.A1(\data_array.data1[12][38] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][38] ),
    .C1(_05066_),
    .X(_05067_));
 sky130_fd_sc_hd__a22o_2 _07865_ (.A1(\data_array.data1[5][38] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][38] ),
    .X(_05068_));
 sky130_fd_sc_hd__a221o_2 _07866_ (.A1(\data_array.data1[4][38] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][38] ),
    .C1(_05068_),
    .X(_05069_));
 sky130_fd_sc_hd__a22o_2 _07867_ (.A1(_03506_),
    .A2(_05063_),
    .B1(_05067_),
    .B2(_03522_),
    .X(_05070_));
 sky130_fd_sc_hd__a22o_2 _07868_ (.A1(_03518_),
    .A2(_05065_),
    .B1(_05069_),
    .B2(_03526_),
    .X(_05071_));
 sky130_fd_sc_hd__or2_2 _07869_ (.A(_05070_),
    .B(_05071_),
    .X(_00095_));
 sky130_fd_sc_hd__a22o_2 _07870_ (.A1(\data_array.data1[9][39] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][39] ),
    .X(_05072_));
 sky130_fd_sc_hd__a221o_2 _07871_ (.A1(\data_array.data1[8][39] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][39] ),
    .C1(_05072_),
    .X(_05073_));
 sky130_fd_sc_hd__a22o_2 _07872_ (.A1(\data_array.data1[1][39] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][39] ),
    .X(_05074_));
 sky130_fd_sc_hd__a221o_2 _07873_ (.A1(\data_array.data1[0][39] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][39] ),
    .C1(_05074_),
    .X(_05075_));
 sky130_fd_sc_hd__a22o_2 _07874_ (.A1(\data_array.data1[13][39] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][39] ),
    .X(_05076_));
 sky130_fd_sc_hd__a221o_2 _07875_ (.A1(\data_array.data1[12][39] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][39] ),
    .C1(_05076_),
    .X(_05077_));
 sky130_fd_sc_hd__a22o_2 _07876_ (.A1(\data_array.data1[5][39] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][39] ),
    .X(_05078_));
 sky130_fd_sc_hd__a221o_2 _07877_ (.A1(\data_array.data1[4][39] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][39] ),
    .C1(_05078_),
    .X(_05079_));
 sky130_fd_sc_hd__a22o_2 _07878_ (.A1(_03506_),
    .A2(_05073_),
    .B1(_05077_),
    .B2(_03522_),
    .X(_05080_));
 sky130_fd_sc_hd__a22o_2 _07879_ (.A1(_03518_),
    .A2(_05075_),
    .B1(_05079_),
    .B2(_03526_),
    .X(_05081_));
 sky130_fd_sc_hd__or2_2 _07880_ (.A(_05080_),
    .B(_05081_),
    .X(_00096_));
 sky130_fd_sc_hd__a22o_2 _07881_ (.A1(\data_array.data1[13][40] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][40] ),
    .X(_05082_));
 sky130_fd_sc_hd__a221o_2 _07882_ (.A1(\data_array.data1[12][40] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][40] ),
    .C1(_05082_),
    .X(_05083_));
 sky130_fd_sc_hd__a22o_2 _07883_ (.A1(\data_array.data1[5][40] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][40] ),
    .X(_05084_));
 sky130_fd_sc_hd__a221o_2 _07884_ (.A1(\data_array.data1[4][40] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][40] ),
    .C1(_05084_),
    .X(_05085_));
 sky130_fd_sc_hd__a22o_2 _07885_ (.A1(\data_array.data1[9][40] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][40] ),
    .X(_05086_));
 sky130_fd_sc_hd__a221o_2 _07886_ (.A1(\data_array.data1[8][40] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][40] ),
    .C1(_05086_),
    .X(_05087_));
 sky130_fd_sc_hd__a22o_2 _07887_ (.A1(\data_array.data1[1][40] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][40] ),
    .X(_05088_));
 sky130_fd_sc_hd__a221o_2 _07888_ (.A1(\data_array.data1[0][40] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][40] ),
    .C1(_05088_),
    .X(_05089_));
 sky130_fd_sc_hd__a22o_2 _07889_ (.A1(_03522_),
    .A2(_05083_),
    .B1(_05087_),
    .B2(_03506_),
    .X(_05090_));
 sky130_fd_sc_hd__a22o_2 _07890_ (.A1(_03526_),
    .A2(_05085_),
    .B1(_05089_),
    .B2(_03518_),
    .X(_05091_));
 sky130_fd_sc_hd__or2_2 _07891_ (.A(_05090_),
    .B(_05091_),
    .X(_00098_));
 sky130_fd_sc_hd__a22o_2 _07892_ (.A1(\data_array.data1[9][41] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][41] ),
    .X(_05092_));
 sky130_fd_sc_hd__a221o_2 _07893_ (.A1(\data_array.data1[8][41] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][41] ),
    .C1(_05092_),
    .X(_05093_));
 sky130_fd_sc_hd__a22o_2 _07894_ (.A1(\data_array.data1[5][41] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][41] ),
    .X(_05094_));
 sky130_fd_sc_hd__a221o_2 _07895_ (.A1(\data_array.data1[4][41] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][41] ),
    .C1(_05094_),
    .X(_05095_));
 sky130_fd_sc_hd__a22o_2 _07896_ (.A1(\data_array.data1[13][41] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][41] ),
    .X(_05096_));
 sky130_fd_sc_hd__a221o_2 _07897_ (.A1(\data_array.data1[12][41] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][41] ),
    .C1(_05096_),
    .X(_05097_));
 sky130_fd_sc_hd__a22o_2 _07898_ (.A1(\data_array.data1[1][41] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][41] ),
    .X(_05098_));
 sky130_fd_sc_hd__a221o_2 _07899_ (.A1(\data_array.data1[0][41] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][41] ),
    .C1(_05098_),
    .X(_05099_));
 sky130_fd_sc_hd__a22o_2 _07900_ (.A1(_03506_),
    .A2(_05093_),
    .B1(_05097_),
    .B2(_03522_),
    .X(_05100_));
 sky130_fd_sc_hd__a22o_2 _07901_ (.A1(_03526_),
    .A2(_05095_),
    .B1(_05099_),
    .B2(_03518_),
    .X(_05101_));
 sky130_fd_sc_hd__or2_2 _07902_ (.A(_05100_),
    .B(_05101_),
    .X(_00099_));
 sky130_fd_sc_hd__a22o_2 _07903_ (.A1(\data_array.data1[9][42] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][42] ),
    .X(_05102_));
 sky130_fd_sc_hd__a221o_2 _07904_ (.A1(\data_array.data1[8][42] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][42] ),
    .C1(_05102_),
    .X(_05103_));
 sky130_fd_sc_hd__a22o_2 _07905_ (.A1(\data_array.data1[5][42] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][42] ),
    .X(_05104_));
 sky130_fd_sc_hd__a221o_2 _07906_ (.A1(\data_array.data1[4][42] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][42] ),
    .C1(_05104_),
    .X(_05105_));
 sky130_fd_sc_hd__a22o_2 _07907_ (.A1(\data_array.data1[13][42] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][42] ),
    .X(_05106_));
 sky130_fd_sc_hd__a221o_2 _07908_ (.A1(\data_array.data1[12][42] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][42] ),
    .C1(_05106_),
    .X(_05107_));
 sky130_fd_sc_hd__a22o_2 _07909_ (.A1(\data_array.data1[1][42] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][42] ),
    .X(_05108_));
 sky130_fd_sc_hd__a221o_2 _07910_ (.A1(\data_array.data1[0][42] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][42] ),
    .C1(_05108_),
    .X(_05109_));
 sky130_fd_sc_hd__a22o_2 _07911_ (.A1(_03506_),
    .A2(_05103_),
    .B1(_05107_),
    .B2(_03522_),
    .X(_05110_));
 sky130_fd_sc_hd__a22o_2 _07912_ (.A1(_03526_),
    .A2(_05105_),
    .B1(_05109_),
    .B2(_03518_),
    .X(_05111_));
 sky130_fd_sc_hd__or2_2 _07913_ (.A(_05110_),
    .B(_05111_),
    .X(_00100_));
 sky130_fd_sc_hd__a22o_2 _07914_ (.A1(\data_array.data1[9][43] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][43] ),
    .X(_05112_));
 sky130_fd_sc_hd__a221o_2 _07915_ (.A1(\data_array.data1[8][43] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][43] ),
    .C1(_05112_),
    .X(_05113_));
 sky130_fd_sc_hd__a22o_2 _07916_ (.A1(\data_array.data1[1][43] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][43] ),
    .X(_05114_));
 sky130_fd_sc_hd__a221o_2 _07917_ (.A1(\data_array.data1[0][43] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][43] ),
    .C1(_05114_),
    .X(_05115_));
 sky130_fd_sc_hd__a22o_2 _07918_ (.A1(\data_array.data1[13][43] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][43] ),
    .X(_05116_));
 sky130_fd_sc_hd__a221o_2 _07919_ (.A1(\data_array.data1[12][43] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][43] ),
    .C1(_05116_),
    .X(_05117_));
 sky130_fd_sc_hd__a22o_2 _07920_ (.A1(\data_array.data1[5][43] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][43] ),
    .X(_05118_));
 sky130_fd_sc_hd__a221o_2 _07921_ (.A1(\data_array.data1[4][43] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][43] ),
    .C1(_05118_),
    .X(_05119_));
 sky130_fd_sc_hd__a22o_2 _07922_ (.A1(_03506_),
    .A2(_05113_),
    .B1(_05117_),
    .B2(_03522_),
    .X(_05120_));
 sky130_fd_sc_hd__a22o_2 _07923_ (.A1(_03518_),
    .A2(_05115_),
    .B1(_05119_),
    .B2(_03526_),
    .X(_05121_));
 sky130_fd_sc_hd__or2_2 _07924_ (.A(_05120_),
    .B(_05121_),
    .X(_00101_));
 sky130_fd_sc_hd__a22o_2 _07925_ (.A1(\data_array.data1[9][44] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][44] ),
    .X(_05122_));
 sky130_fd_sc_hd__a221o_2 _07926_ (.A1(\data_array.data1[8][44] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][44] ),
    .C1(_05122_),
    .X(_05123_));
 sky130_fd_sc_hd__a22o_2 _07927_ (.A1(\data_array.data1[1][44] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][44] ),
    .X(_05124_));
 sky130_fd_sc_hd__a221o_2 _07928_ (.A1(\data_array.data1[0][44] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][44] ),
    .C1(_05124_),
    .X(_05125_));
 sky130_fd_sc_hd__a22o_2 _07929_ (.A1(\data_array.data1[13][44] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][44] ),
    .X(_05126_));
 sky130_fd_sc_hd__a221o_2 _07930_ (.A1(\data_array.data1[12][44] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][44] ),
    .C1(_05126_),
    .X(_05127_));
 sky130_fd_sc_hd__a22o_2 _07931_ (.A1(\data_array.data1[5][44] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][44] ),
    .X(_05128_));
 sky130_fd_sc_hd__a221o_2 _07932_ (.A1(\data_array.data1[4][44] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][44] ),
    .C1(_05128_),
    .X(_05129_));
 sky130_fd_sc_hd__a22o_2 _07933_ (.A1(_03506_),
    .A2(_05123_),
    .B1(_05127_),
    .B2(_03522_),
    .X(_05130_));
 sky130_fd_sc_hd__a22o_2 _07934_ (.A1(_03518_),
    .A2(_05125_),
    .B1(_05129_),
    .B2(_03526_),
    .X(_05131_));
 sky130_fd_sc_hd__or2_2 _07935_ (.A(_05130_),
    .B(_05131_),
    .X(_00102_));
 sky130_fd_sc_hd__a22o_2 _07936_ (.A1(\data_array.data1[13][45] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][45] ),
    .X(_05132_));
 sky130_fd_sc_hd__a221o_2 _07937_ (.A1(\data_array.data1[12][45] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][45] ),
    .C1(_05132_),
    .X(_05133_));
 sky130_fd_sc_hd__a22o_2 _07938_ (.A1(\data_array.data1[1][45] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][45] ),
    .X(_05134_));
 sky130_fd_sc_hd__a221o_2 _07939_ (.A1(\data_array.data1[0][45] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][45] ),
    .C1(_05134_),
    .X(_05135_));
 sky130_fd_sc_hd__a22o_2 _07940_ (.A1(\data_array.data1[9][45] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][45] ),
    .X(_05136_));
 sky130_fd_sc_hd__a221o_2 _07941_ (.A1(\data_array.data1[8][45] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][45] ),
    .C1(_05136_),
    .X(_05137_));
 sky130_fd_sc_hd__a22o_2 _07942_ (.A1(\data_array.data1[5][45] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][45] ),
    .X(_05138_));
 sky130_fd_sc_hd__a221o_2 _07943_ (.A1(\data_array.data1[4][45] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][45] ),
    .C1(_05138_),
    .X(_05139_));
 sky130_fd_sc_hd__a22o_2 _07944_ (.A1(_03522_),
    .A2(_05133_),
    .B1(_05137_),
    .B2(_03506_),
    .X(_05140_));
 sky130_fd_sc_hd__a22o_2 _07945_ (.A1(_03518_),
    .A2(_05135_),
    .B1(_05139_),
    .B2(_03526_),
    .X(_05141_));
 sky130_fd_sc_hd__or2_2 _07946_ (.A(_05140_),
    .B(_05141_),
    .X(_00103_));
 sky130_fd_sc_hd__a22o_2 _07947_ (.A1(\data_array.data1[9][46] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][46] ),
    .X(_05142_));
 sky130_fd_sc_hd__a221o_2 _07948_ (.A1(\data_array.data1[8][46] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][46] ),
    .C1(_05142_),
    .X(_05143_));
 sky130_fd_sc_hd__a22o_2 _07949_ (.A1(\data_array.data1[5][46] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][46] ),
    .X(_05144_));
 sky130_fd_sc_hd__a221o_2 _07950_ (.A1(\data_array.data1[4][46] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][46] ),
    .C1(_05144_),
    .X(_05145_));
 sky130_fd_sc_hd__a22o_2 _07951_ (.A1(\data_array.data1[13][46] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][46] ),
    .X(_05146_));
 sky130_fd_sc_hd__a221o_2 _07952_ (.A1(\data_array.data1[12][46] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][46] ),
    .C1(_05146_),
    .X(_05147_));
 sky130_fd_sc_hd__a22o_2 _07953_ (.A1(\data_array.data1[1][46] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][46] ),
    .X(_05148_));
 sky130_fd_sc_hd__a221o_2 _07954_ (.A1(\data_array.data1[0][46] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][46] ),
    .C1(_05148_),
    .X(_05149_));
 sky130_fd_sc_hd__a22o_2 _07955_ (.A1(_03506_),
    .A2(_05143_),
    .B1(_05147_),
    .B2(_03522_),
    .X(_05150_));
 sky130_fd_sc_hd__a22o_2 _07956_ (.A1(_03526_),
    .A2(_05145_),
    .B1(_05149_),
    .B2(_03518_),
    .X(_05151_));
 sky130_fd_sc_hd__or2_2 _07957_ (.A(_05150_),
    .B(_05151_),
    .X(_00104_));
 sky130_fd_sc_hd__a22o_2 _07958_ (.A1(\data_array.data1[9][47] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][47] ),
    .X(_05152_));
 sky130_fd_sc_hd__a221o_2 _07959_ (.A1(\data_array.data1[8][47] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][47] ),
    .C1(_05152_),
    .X(_05153_));
 sky130_fd_sc_hd__a22o_2 _07960_ (.A1(\data_array.data1[5][47] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][47] ),
    .X(_05154_));
 sky130_fd_sc_hd__a221o_2 _07961_ (.A1(\data_array.data1[4][47] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][47] ),
    .C1(_05154_),
    .X(_05155_));
 sky130_fd_sc_hd__a22o_2 _07962_ (.A1(\data_array.data1[13][47] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][47] ),
    .X(_05156_));
 sky130_fd_sc_hd__a221o_2 _07963_ (.A1(\data_array.data1[12][47] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][47] ),
    .C1(_05156_),
    .X(_05157_));
 sky130_fd_sc_hd__a22o_2 _07964_ (.A1(\data_array.data1[1][47] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][47] ),
    .X(_05158_));
 sky130_fd_sc_hd__a221o_2 _07965_ (.A1(\data_array.data1[0][47] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][47] ),
    .C1(_05158_),
    .X(_05159_));
 sky130_fd_sc_hd__a22o_2 _07966_ (.A1(_03506_),
    .A2(_05153_),
    .B1(_05157_),
    .B2(_03522_),
    .X(_05160_));
 sky130_fd_sc_hd__a22o_2 _07967_ (.A1(_03526_),
    .A2(_05155_),
    .B1(_05159_),
    .B2(_03518_),
    .X(_05161_));
 sky130_fd_sc_hd__or2_2 _07968_ (.A(_05160_),
    .B(_05161_),
    .X(_00105_));
 sky130_fd_sc_hd__a22o_2 _07969_ (.A1(\data_array.data1[9][48] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][48] ),
    .X(_05162_));
 sky130_fd_sc_hd__a221o_2 _07970_ (.A1(\data_array.data1[8][48] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][48] ),
    .C1(_05162_),
    .X(_05163_));
 sky130_fd_sc_hd__a22o_2 _07971_ (.A1(\data_array.data1[5][48] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][48] ),
    .X(_05164_));
 sky130_fd_sc_hd__a221o_2 _07972_ (.A1(\data_array.data1[4][48] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][48] ),
    .C1(_05164_),
    .X(_05165_));
 sky130_fd_sc_hd__a22o_2 _07973_ (.A1(\data_array.data1[13][48] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][48] ),
    .X(_05166_));
 sky130_fd_sc_hd__a221o_2 _07974_ (.A1(\data_array.data1[12][48] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][48] ),
    .C1(_05166_),
    .X(_05167_));
 sky130_fd_sc_hd__a22o_2 _07975_ (.A1(\data_array.data1[1][48] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][48] ),
    .X(_05168_));
 sky130_fd_sc_hd__a221o_2 _07976_ (.A1(\data_array.data1[0][48] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][48] ),
    .C1(_05168_),
    .X(_05169_));
 sky130_fd_sc_hd__a22o_2 _07977_ (.A1(_03506_),
    .A2(_05163_),
    .B1(_05167_),
    .B2(_03522_),
    .X(_05170_));
 sky130_fd_sc_hd__a22o_2 _07978_ (.A1(_03526_),
    .A2(_05165_),
    .B1(_05169_),
    .B2(_03518_),
    .X(_05171_));
 sky130_fd_sc_hd__or2_2 _07979_ (.A(_05170_),
    .B(_05171_),
    .X(_00106_));
 sky130_fd_sc_hd__a22o_2 _07980_ (.A1(\data_array.data1[13][49] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][49] ),
    .X(_05172_));
 sky130_fd_sc_hd__a221o_2 _07981_ (.A1(\data_array.data1[12][49] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][49] ),
    .C1(_05172_),
    .X(_05173_));
 sky130_fd_sc_hd__a22o_2 _07982_ (.A1(\data_array.data1[1][49] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][49] ),
    .X(_05174_));
 sky130_fd_sc_hd__a221o_2 _07983_ (.A1(\data_array.data1[0][49] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][49] ),
    .C1(_05174_),
    .X(_05175_));
 sky130_fd_sc_hd__a22o_2 _07984_ (.A1(\data_array.data1[9][49] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][49] ),
    .X(_05176_));
 sky130_fd_sc_hd__a221o_2 _07985_ (.A1(\data_array.data1[8][49] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][49] ),
    .C1(_05176_),
    .X(_05177_));
 sky130_fd_sc_hd__a22o_2 _07986_ (.A1(\data_array.data1[5][49] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][49] ),
    .X(_05178_));
 sky130_fd_sc_hd__a221o_2 _07987_ (.A1(\data_array.data1[4][49] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][49] ),
    .C1(_05178_),
    .X(_05179_));
 sky130_fd_sc_hd__a22o_2 _07988_ (.A1(_03522_),
    .A2(_05173_),
    .B1(_05177_),
    .B2(_03506_),
    .X(_05180_));
 sky130_fd_sc_hd__a22o_2 _07989_ (.A1(_03518_),
    .A2(_05175_),
    .B1(_05179_),
    .B2(_03526_),
    .X(_05181_));
 sky130_fd_sc_hd__or2_2 _07990_ (.A(_05180_),
    .B(_05181_),
    .X(_00107_));
 sky130_fd_sc_hd__a22o_2 _07991_ (.A1(\data_array.data1[9][50] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][50] ),
    .X(_05182_));
 sky130_fd_sc_hd__a221o_2 _07992_ (.A1(\data_array.data1[8][50] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][50] ),
    .C1(_05182_),
    .X(_05183_));
 sky130_fd_sc_hd__a22o_2 _07993_ (.A1(\data_array.data1[5][50] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][50] ),
    .X(_05184_));
 sky130_fd_sc_hd__a221o_2 _07994_ (.A1(\data_array.data1[4][50] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][50] ),
    .C1(_05184_),
    .X(_05185_));
 sky130_fd_sc_hd__a22o_2 _07995_ (.A1(\data_array.data1[13][50] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][50] ),
    .X(_05186_));
 sky130_fd_sc_hd__a221o_2 _07996_ (.A1(\data_array.data1[12][50] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][50] ),
    .C1(_05186_),
    .X(_05187_));
 sky130_fd_sc_hd__a22o_2 _07997_ (.A1(\data_array.data1[1][50] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][50] ),
    .X(_05188_));
 sky130_fd_sc_hd__a221o_2 _07998_ (.A1(\data_array.data1[0][50] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][50] ),
    .C1(_05188_),
    .X(_05189_));
 sky130_fd_sc_hd__a22o_2 _07999_ (.A1(_03506_),
    .A2(_05183_),
    .B1(_05187_),
    .B2(_03522_),
    .X(_05190_));
 sky130_fd_sc_hd__a22o_2 _08000_ (.A1(_03526_),
    .A2(_05185_),
    .B1(_05189_),
    .B2(_03518_),
    .X(_05191_));
 sky130_fd_sc_hd__or2_2 _08001_ (.A(_05190_),
    .B(_05191_),
    .X(_00109_));
 sky130_fd_sc_hd__a22o_2 _08002_ (.A1(\data_array.data1[13][51] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][51] ),
    .X(_05192_));
 sky130_fd_sc_hd__a221o_2 _08003_ (.A1(\data_array.data1[12][51] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][51] ),
    .C1(_05192_),
    .X(_05193_));
 sky130_fd_sc_hd__a22o_2 _08004_ (.A1(\data_array.data1[5][51] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][51] ),
    .X(_05194_));
 sky130_fd_sc_hd__a221o_2 _08005_ (.A1(\data_array.data1[4][51] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][51] ),
    .C1(_05194_),
    .X(_05195_));
 sky130_fd_sc_hd__a22o_2 _08006_ (.A1(\data_array.data1[9][51] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][51] ),
    .X(_05196_));
 sky130_fd_sc_hd__a221o_2 _08007_ (.A1(\data_array.data1[8][51] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][51] ),
    .C1(_05196_),
    .X(_05197_));
 sky130_fd_sc_hd__a22o_2 _08008_ (.A1(\data_array.data1[1][51] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][51] ),
    .X(_05198_));
 sky130_fd_sc_hd__a221o_2 _08009_ (.A1(\data_array.data1[0][51] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][51] ),
    .C1(_05198_),
    .X(_05199_));
 sky130_fd_sc_hd__a22o_2 _08010_ (.A1(_03522_),
    .A2(_05193_),
    .B1(_05197_),
    .B2(_03506_),
    .X(_05200_));
 sky130_fd_sc_hd__a22o_2 _08011_ (.A1(_03526_),
    .A2(_05195_),
    .B1(_05199_),
    .B2(_03518_),
    .X(_05201_));
 sky130_fd_sc_hd__or2_2 _08012_ (.A(_05200_),
    .B(_05201_),
    .X(_00110_));
 sky130_fd_sc_hd__a22o_2 _08013_ (.A1(\data_array.data1[13][52] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][52] ),
    .X(_05202_));
 sky130_fd_sc_hd__a221o_2 _08014_ (.A1(\data_array.data1[12][52] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][52] ),
    .C1(_05202_),
    .X(_05203_));
 sky130_fd_sc_hd__a22o_2 _08015_ (.A1(\data_array.data1[5][52] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][52] ),
    .X(_05204_));
 sky130_fd_sc_hd__a221o_2 _08016_ (.A1(\data_array.data1[4][52] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][52] ),
    .C1(_05204_),
    .X(_05205_));
 sky130_fd_sc_hd__a22o_2 _08017_ (.A1(\data_array.data1[9][52] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][52] ),
    .X(_05206_));
 sky130_fd_sc_hd__a221o_2 _08018_ (.A1(\data_array.data1[8][52] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][52] ),
    .C1(_05206_),
    .X(_05207_));
 sky130_fd_sc_hd__a22o_2 _08019_ (.A1(\data_array.data1[1][52] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][52] ),
    .X(_05208_));
 sky130_fd_sc_hd__a221o_2 _08020_ (.A1(\data_array.data1[0][52] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][52] ),
    .C1(_05208_),
    .X(_05209_));
 sky130_fd_sc_hd__a22o_2 _08021_ (.A1(_03522_),
    .A2(_05203_),
    .B1(_05207_),
    .B2(_03506_),
    .X(_05210_));
 sky130_fd_sc_hd__a22o_2 _08022_ (.A1(_03526_),
    .A2(_05205_),
    .B1(_05209_),
    .B2(_03518_),
    .X(_05211_));
 sky130_fd_sc_hd__or2_2 _08023_ (.A(_05210_),
    .B(_05211_),
    .X(_00111_));
 sky130_fd_sc_hd__a22o_2 _08024_ (.A1(\data_array.data1[9][53] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][53] ),
    .X(_05212_));
 sky130_fd_sc_hd__a221o_2 _08025_ (.A1(\data_array.data1[8][53] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][53] ),
    .C1(_05212_),
    .X(_05213_));
 sky130_fd_sc_hd__a22o_2 _08026_ (.A1(\data_array.data1[1][53] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][53] ),
    .X(_05214_));
 sky130_fd_sc_hd__a221o_2 _08027_ (.A1(\data_array.data1[0][53] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][53] ),
    .C1(_05214_),
    .X(_05215_));
 sky130_fd_sc_hd__a22o_2 _08028_ (.A1(\data_array.data1[13][53] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][53] ),
    .X(_05216_));
 sky130_fd_sc_hd__a221o_2 _08029_ (.A1(\data_array.data1[12][53] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][53] ),
    .C1(_05216_),
    .X(_05217_));
 sky130_fd_sc_hd__a22o_2 _08030_ (.A1(\data_array.data1[5][53] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][53] ),
    .X(_05218_));
 sky130_fd_sc_hd__a221o_2 _08031_ (.A1(\data_array.data1[4][53] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][53] ),
    .C1(_05218_),
    .X(_05219_));
 sky130_fd_sc_hd__a22o_2 _08032_ (.A1(_03506_),
    .A2(_05213_),
    .B1(_05217_),
    .B2(_03522_),
    .X(_05220_));
 sky130_fd_sc_hd__a22o_2 _08033_ (.A1(_03518_),
    .A2(_05215_),
    .B1(_05219_),
    .B2(_03526_),
    .X(_05221_));
 sky130_fd_sc_hd__or2_2 _08034_ (.A(_05220_),
    .B(_05221_),
    .X(_00112_));
 sky130_fd_sc_hd__a22o_2 _08035_ (.A1(\data_array.data1[9][54] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][54] ),
    .X(_05222_));
 sky130_fd_sc_hd__a221o_2 _08036_ (.A1(\data_array.data1[8][54] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][54] ),
    .C1(_05222_),
    .X(_05223_));
 sky130_fd_sc_hd__a22o_2 _08037_ (.A1(\data_array.data1[1][54] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][54] ),
    .X(_05224_));
 sky130_fd_sc_hd__a221o_2 _08038_ (.A1(\data_array.data1[0][54] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][54] ),
    .C1(_05224_),
    .X(_05225_));
 sky130_fd_sc_hd__a22o_2 _08039_ (.A1(\data_array.data1[13][54] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][54] ),
    .X(_05226_));
 sky130_fd_sc_hd__a221o_2 _08040_ (.A1(\data_array.data1[12][54] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][54] ),
    .C1(_05226_),
    .X(_05227_));
 sky130_fd_sc_hd__a22o_2 _08041_ (.A1(\data_array.data1[5][54] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][54] ),
    .X(_05228_));
 sky130_fd_sc_hd__a221o_2 _08042_ (.A1(\data_array.data1[4][54] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][54] ),
    .C1(_05228_),
    .X(_05229_));
 sky130_fd_sc_hd__a22o_2 _08043_ (.A1(_03506_),
    .A2(_05223_),
    .B1(_05227_),
    .B2(_03522_),
    .X(_05230_));
 sky130_fd_sc_hd__a22o_2 _08044_ (.A1(_03518_),
    .A2(_05225_),
    .B1(_05229_),
    .B2(_03526_),
    .X(_05231_));
 sky130_fd_sc_hd__or2_2 _08045_ (.A(_05230_),
    .B(_05231_),
    .X(_00113_));
 sky130_fd_sc_hd__a22o_2 _08046_ (.A1(\data_array.data1[13][55] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][55] ),
    .X(_05232_));
 sky130_fd_sc_hd__a221o_2 _08047_ (.A1(\data_array.data1[12][55] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][55] ),
    .C1(_05232_),
    .X(_05233_));
 sky130_fd_sc_hd__a22o_2 _08048_ (.A1(\data_array.data1[1][55] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][55] ),
    .X(_05234_));
 sky130_fd_sc_hd__a221o_2 _08049_ (.A1(\data_array.data1[0][55] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][55] ),
    .C1(_05234_),
    .X(_05235_));
 sky130_fd_sc_hd__a22o_2 _08050_ (.A1(\data_array.data1[9][55] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][55] ),
    .X(_05236_));
 sky130_fd_sc_hd__a221o_2 _08051_ (.A1(\data_array.data1[8][55] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][55] ),
    .C1(_05236_),
    .X(_05237_));
 sky130_fd_sc_hd__a22o_2 _08052_ (.A1(\data_array.data1[5][55] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][55] ),
    .X(_05238_));
 sky130_fd_sc_hd__a221o_2 _08053_ (.A1(\data_array.data1[4][55] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][55] ),
    .C1(_05238_),
    .X(_05239_));
 sky130_fd_sc_hd__a22o_2 _08054_ (.A1(_03522_),
    .A2(_05233_),
    .B1(_05237_),
    .B2(_03506_),
    .X(_05240_));
 sky130_fd_sc_hd__a22o_2 _08055_ (.A1(_03518_),
    .A2(_05235_),
    .B1(_05239_),
    .B2(_03526_),
    .X(_05241_));
 sky130_fd_sc_hd__or2_2 _08056_ (.A(_05240_),
    .B(_05241_),
    .X(_00114_));
 sky130_fd_sc_hd__a22o_2 _08057_ (.A1(\data_array.data1[13][56] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][56] ),
    .X(_05242_));
 sky130_fd_sc_hd__a221o_2 _08058_ (.A1(\data_array.data1[12][56] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][56] ),
    .C1(_05242_),
    .X(_05243_));
 sky130_fd_sc_hd__a22o_2 _08059_ (.A1(\data_array.data1[5][56] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][56] ),
    .X(_05244_));
 sky130_fd_sc_hd__a221o_2 _08060_ (.A1(\data_array.data1[4][56] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][56] ),
    .C1(_05244_),
    .X(_05245_));
 sky130_fd_sc_hd__a22o_2 _08061_ (.A1(\data_array.data1[9][56] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][56] ),
    .X(_05246_));
 sky130_fd_sc_hd__a221o_2 _08062_ (.A1(\data_array.data1[8][56] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][56] ),
    .C1(_05246_),
    .X(_05247_));
 sky130_fd_sc_hd__a22o_2 _08063_ (.A1(\data_array.data1[1][56] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][56] ),
    .X(_05248_));
 sky130_fd_sc_hd__a221o_2 _08064_ (.A1(\data_array.data1[0][56] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][56] ),
    .C1(_05248_),
    .X(_05249_));
 sky130_fd_sc_hd__a22o_2 _08065_ (.A1(_03522_),
    .A2(_05243_),
    .B1(_05247_),
    .B2(_03506_),
    .X(_05250_));
 sky130_fd_sc_hd__a22o_2 _08066_ (.A1(_03526_),
    .A2(_05245_),
    .B1(_05249_),
    .B2(_03518_),
    .X(_05251_));
 sky130_fd_sc_hd__or2_2 _08067_ (.A(_05250_),
    .B(_05251_),
    .X(_00115_));
 sky130_fd_sc_hd__a22o_2 _08068_ (.A1(\data_array.data1[13][57] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][57] ),
    .X(_05252_));
 sky130_fd_sc_hd__a221o_2 _08069_ (.A1(\data_array.data1[12][57] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][57] ),
    .C1(_05252_),
    .X(_05253_));
 sky130_fd_sc_hd__a22o_2 _08070_ (.A1(\data_array.data1[1][57] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][57] ),
    .X(_05254_));
 sky130_fd_sc_hd__a221o_2 _08071_ (.A1(\data_array.data1[0][57] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][57] ),
    .C1(_05254_),
    .X(_05255_));
 sky130_fd_sc_hd__a22o_2 _08072_ (.A1(\data_array.data1[9][57] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][57] ),
    .X(_05256_));
 sky130_fd_sc_hd__a221o_2 _08073_ (.A1(\data_array.data1[8][57] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][57] ),
    .C1(_05256_),
    .X(_05257_));
 sky130_fd_sc_hd__a22o_2 _08074_ (.A1(\data_array.data1[5][57] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][57] ),
    .X(_05258_));
 sky130_fd_sc_hd__a221o_2 _08075_ (.A1(\data_array.data1[4][57] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][57] ),
    .C1(_05258_),
    .X(_05259_));
 sky130_fd_sc_hd__a22o_2 _08076_ (.A1(_03522_),
    .A2(_05253_),
    .B1(_05257_),
    .B2(_03506_),
    .X(_05260_));
 sky130_fd_sc_hd__a22o_2 _08077_ (.A1(_03518_),
    .A2(_05255_),
    .B1(_05259_),
    .B2(_03526_),
    .X(_05261_));
 sky130_fd_sc_hd__or2_2 _08078_ (.A(_05260_),
    .B(_05261_),
    .X(_00116_));
 sky130_fd_sc_hd__a22o_2 _08079_ (.A1(\data_array.data1[9][58] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][58] ),
    .X(_05262_));
 sky130_fd_sc_hd__a221o_2 _08080_ (.A1(\data_array.data1[8][58] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][58] ),
    .C1(_05262_),
    .X(_05263_));
 sky130_fd_sc_hd__a22o_2 _08081_ (.A1(\data_array.data1[5][58] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][58] ),
    .X(_05264_));
 sky130_fd_sc_hd__a221o_2 _08082_ (.A1(\data_array.data1[4][58] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][58] ),
    .C1(_05264_),
    .X(_05265_));
 sky130_fd_sc_hd__a22o_2 _08083_ (.A1(\data_array.data1[13][58] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][58] ),
    .X(_05266_));
 sky130_fd_sc_hd__a221o_2 _08084_ (.A1(\data_array.data1[12][58] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][58] ),
    .C1(_05266_),
    .X(_05267_));
 sky130_fd_sc_hd__a22o_2 _08085_ (.A1(\data_array.data1[1][58] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][58] ),
    .X(_05268_));
 sky130_fd_sc_hd__a221o_2 _08086_ (.A1(\data_array.data1[0][58] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][58] ),
    .C1(_05268_),
    .X(_05269_));
 sky130_fd_sc_hd__a22o_2 _08087_ (.A1(_03506_),
    .A2(_05263_),
    .B1(_05267_),
    .B2(_03522_),
    .X(_05270_));
 sky130_fd_sc_hd__a22o_2 _08088_ (.A1(_03526_),
    .A2(_05265_),
    .B1(_05269_),
    .B2(_03518_),
    .X(_05271_));
 sky130_fd_sc_hd__or2_2 _08089_ (.A(_05270_),
    .B(_05271_),
    .X(_00117_));
 sky130_fd_sc_hd__a22o_2 _08090_ (.A1(\data_array.data1[9][59] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][59] ),
    .X(_05272_));
 sky130_fd_sc_hd__a221o_2 _08091_ (.A1(\data_array.data1[8][59] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][59] ),
    .C1(_05272_),
    .X(_05273_));
 sky130_fd_sc_hd__a22o_2 _08092_ (.A1(\data_array.data1[1][59] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][59] ),
    .X(_05274_));
 sky130_fd_sc_hd__a221o_2 _08093_ (.A1(\data_array.data1[0][59] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][59] ),
    .C1(_05274_),
    .X(_05275_));
 sky130_fd_sc_hd__a22o_2 _08094_ (.A1(\data_array.data1[13][59] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][59] ),
    .X(_05276_));
 sky130_fd_sc_hd__a221o_2 _08095_ (.A1(\data_array.data1[12][59] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][59] ),
    .C1(_05276_),
    .X(_05277_));
 sky130_fd_sc_hd__a22o_2 _08096_ (.A1(\data_array.data1[5][59] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][59] ),
    .X(_05278_));
 sky130_fd_sc_hd__a221o_2 _08097_ (.A1(\data_array.data1[4][59] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][59] ),
    .C1(_05278_),
    .X(_05279_));
 sky130_fd_sc_hd__a22o_2 _08098_ (.A1(_03506_),
    .A2(_05273_),
    .B1(_05277_),
    .B2(_03522_),
    .X(_05280_));
 sky130_fd_sc_hd__a22o_2 _08099_ (.A1(_03518_),
    .A2(_05275_),
    .B1(_05279_),
    .B2(_03526_),
    .X(_05281_));
 sky130_fd_sc_hd__or2_2 _08100_ (.A(_05280_),
    .B(_05281_),
    .X(_00118_));
 sky130_fd_sc_hd__a22o_2 _08101_ (.A1(\data_array.data1[9][60] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][60] ),
    .X(_05282_));
 sky130_fd_sc_hd__a221o_2 _08102_ (.A1(\data_array.data1[8][60] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][60] ),
    .C1(_05282_),
    .X(_05283_));
 sky130_fd_sc_hd__a22o_2 _08103_ (.A1(\data_array.data1[5][60] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][60] ),
    .X(_05284_));
 sky130_fd_sc_hd__a221o_2 _08104_ (.A1(\data_array.data1[4][60] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][60] ),
    .C1(_05284_),
    .X(_05285_));
 sky130_fd_sc_hd__a22o_2 _08105_ (.A1(\data_array.data1[13][60] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][60] ),
    .X(_05286_));
 sky130_fd_sc_hd__a221o_2 _08106_ (.A1(\data_array.data1[12][60] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][60] ),
    .C1(_05286_),
    .X(_05287_));
 sky130_fd_sc_hd__a22o_2 _08107_ (.A1(\data_array.data1[1][60] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][60] ),
    .X(_05288_));
 sky130_fd_sc_hd__a221o_2 _08108_ (.A1(\data_array.data1[0][60] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][60] ),
    .C1(_05288_),
    .X(_05289_));
 sky130_fd_sc_hd__a22o_2 _08109_ (.A1(_03506_),
    .A2(_05283_),
    .B1(_05287_),
    .B2(_03522_),
    .X(_05290_));
 sky130_fd_sc_hd__a22o_2 _08110_ (.A1(_03526_),
    .A2(_05285_),
    .B1(_05289_),
    .B2(_03518_),
    .X(_05291_));
 sky130_fd_sc_hd__or2_2 _08111_ (.A(_05290_),
    .B(_05291_),
    .X(_00120_));
 sky130_fd_sc_hd__a22o_2 _08112_ (.A1(\data_array.data1[13][61] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][61] ),
    .X(_05292_));
 sky130_fd_sc_hd__a221o_2 _08113_ (.A1(\data_array.data1[12][61] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][61] ),
    .C1(_05292_),
    .X(_05293_));
 sky130_fd_sc_hd__a22o_2 _08114_ (.A1(\data_array.data1[1][61] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][61] ),
    .X(_05294_));
 sky130_fd_sc_hd__a221o_2 _08115_ (.A1(\data_array.data1[0][61] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][61] ),
    .C1(_05294_),
    .X(_05295_));
 sky130_fd_sc_hd__a22o_2 _08116_ (.A1(\data_array.data1[9][61] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][61] ),
    .X(_05296_));
 sky130_fd_sc_hd__a221o_2 _08117_ (.A1(\data_array.data1[8][61] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][61] ),
    .C1(_05296_),
    .X(_05297_));
 sky130_fd_sc_hd__a22o_2 _08118_ (.A1(\data_array.data1[5][61] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][61] ),
    .X(_05298_));
 sky130_fd_sc_hd__a221o_2 _08119_ (.A1(\data_array.data1[4][61] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][61] ),
    .C1(_05298_),
    .X(_05299_));
 sky130_fd_sc_hd__a22o_2 _08120_ (.A1(_03522_),
    .A2(_05293_),
    .B1(_05297_),
    .B2(_03506_),
    .X(_05300_));
 sky130_fd_sc_hd__a22o_2 _08121_ (.A1(_03518_),
    .A2(_05295_),
    .B1(_05299_),
    .B2(_03526_),
    .X(_05301_));
 sky130_fd_sc_hd__or2_2 _08122_ (.A(_05300_),
    .B(_05301_),
    .X(_00121_));
 sky130_fd_sc_hd__a22o_2 _08123_ (.A1(\data_array.data1[9][62] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][62] ),
    .X(_05302_));
 sky130_fd_sc_hd__a221o_2 _08124_ (.A1(\data_array.data1[8][62] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][62] ),
    .C1(_05302_),
    .X(_05303_));
 sky130_fd_sc_hd__a22o_2 _08125_ (.A1(\data_array.data1[5][62] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][62] ),
    .X(_05304_));
 sky130_fd_sc_hd__a221o_2 _08126_ (.A1(\data_array.data1[4][62] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][62] ),
    .C1(_05304_),
    .X(_05305_));
 sky130_fd_sc_hd__a22o_2 _08127_ (.A1(\data_array.data1[13][62] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][62] ),
    .X(_05306_));
 sky130_fd_sc_hd__a221o_2 _08128_ (.A1(\data_array.data1[12][62] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][62] ),
    .C1(_05306_),
    .X(_05307_));
 sky130_fd_sc_hd__a22o_2 _08129_ (.A1(\data_array.data1[1][62] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][62] ),
    .X(_05308_));
 sky130_fd_sc_hd__a221o_2 _08130_ (.A1(\data_array.data1[0][62] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][62] ),
    .C1(_05308_),
    .X(_05309_));
 sky130_fd_sc_hd__a22o_2 _08131_ (.A1(_03506_),
    .A2(_05303_),
    .B1(_05307_),
    .B2(_03522_),
    .X(_05310_));
 sky130_fd_sc_hd__a22o_2 _08132_ (.A1(_03526_),
    .A2(_05305_),
    .B1(_05309_),
    .B2(_03518_),
    .X(_05311_));
 sky130_fd_sc_hd__or2_2 _08133_ (.A(_05310_),
    .B(_05311_),
    .X(_00122_));
 sky130_fd_sc_hd__a22o_2 _08134_ (.A1(\data_array.data1[13][63] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[14][63] ),
    .X(_05312_));
 sky130_fd_sc_hd__a221o_2 _08135_ (.A1(\data_array.data1[12][63] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[15][63] ),
    .C1(_05312_),
    .X(_05313_));
 sky130_fd_sc_hd__a22o_2 _08136_ (.A1(\data_array.data1[5][63] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[6][63] ),
    .X(_05314_));
 sky130_fd_sc_hd__a221o_2 _08137_ (.A1(\data_array.data1[4][63] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[7][63] ),
    .C1(_05314_),
    .X(_05315_));
 sky130_fd_sc_hd__a22o_2 _08138_ (.A1(\data_array.data1[9][63] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[10][63] ),
    .X(_05316_));
 sky130_fd_sc_hd__a221o_2 _08139_ (.A1(\data_array.data1[8][63] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[11][63] ),
    .C1(_05316_),
    .X(_05317_));
 sky130_fd_sc_hd__a22o_2 _08140_ (.A1(\data_array.data1[1][63] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\data_array.data1[2][63] ),
    .X(_05318_));
 sky130_fd_sc_hd__a221o_2 _08141_ (.A1(\data_array.data1[0][63] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\data_array.data1[3][63] ),
    .C1(_05318_),
    .X(_05319_));
 sky130_fd_sc_hd__a22o_2 _08142_ (.A1(_03522_),
    .A2(_05313_),
    .B1(_05317_),
    .B2(_03506_),
    .X(_05320_));
 sky130_fd_sc_hd__a22o_2 _08143_ (.A1(_03526_),
    .A2(_05315_),
    .B1(_05319_),
    .B2(_03518_),
    .X(_05321_));
 sky130_fd_sc_hd__or2_2 _08144_ (.A(_05320_),
    .B(_05321_),
    .X(_00123_));
 sky130_fd_sc_hd__a22o_2 _08145_ (.A1(\tag_array.dirty1[13] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.dirty1[14] ),
    .X(_05322_));
 sky130_fd_sc_hd__a221o_2 _08146_ (.A1(\tag_array.dirty1[12] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.dirty1[15] ),
    .C1(_05322_),
    .X(_05323_));
 sky130_fd_sc_hd__a22o_2 _08147_ (.A1(\tag_array.dirty1[1] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.dirty1[2] ),
    .X(_05324_));
 sky130_fd_sc_hd__a221o_2 _08148_ (.A1(\tag_array.dirty1[0] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.dirty1[3] ),
    .C1(_05324_),
    .X(_05325_));
 sky130_fd_sc_hd__a22o_2 _08149_ (.A1(\tag_array.dirty1[9] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.dirty1[10] ),
    .X(_05326_));
 sky130_fd_sc_hd__a221o_2 _08150_ (.A1(\tag_array.dirty1[8] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.dirty1[11] ),
    .C1(_05326_),
    .X(_05327_));
 sky130_fd_sc_hd__a22o_2 _08151_ (.A1(\tag_array.dirty1[5] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.dirty1[6] ),
    .X(_05328_));
 sky130_fd_sc_hd__a221o_2 _08152_ (.A1(\tag_array.dirty1[4] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.dirty1[7] ),
    .C1(_05328_),
    .X(_05329_));
 sky130_fd_sc_hd__a22o_2 _08153_ (.A1(_03522_),
    .A2(_05323_),
    .B1(_05327_),
    .B2(_03506_),
    .X(_05330_));
 sky130_fd_sc_hd__a22o_2 _08154_ (.A1(_03518_),
    .A2(_05325_),
    .B1(_05329_),
    .B2(_03526_),
    .X(_05331_));
 sky130_fd_sc_hd__or2_2 _08155_ (.A(_05330_),
    .B(_05331_),
    .X(_00130_));
 sky130_fd_sc_hd__a22o_2 _08156_ (.A1(\tag_array.dirty0[13] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.dirty0[14] ),
    .X(_05332_));
 sky130_fd_sc_hd__a221o_2 _08157_ (.A1(\tag_array.dirty0[12] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.dirty0[15] ),
    .C1(_05332_),
    .X(_05333_));
 sky130_fd_sc_hd__a22o_2 _08158_ (.A1(\tag_array.dirty0[1] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.dirty0[2] ),
    .X(_05334_));
 sky130_fd_sc_hd__a221o_2 _08159_ (.A1(\tag_array.dirty0[0] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.dirty0[3] ),
    .C1(_05334_),
    .X(_05335_));
 sky130_fd_sc_hd__a22o_2 _08160_ (.A1(\tag_array.dirty0[9] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.dirty0[10] ),
    .X(_05336_));
 sky130_fd_sc_hd__a221o_2 _08161_ (.A1(\tag_array.dirty0[8] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.dirty0[11] ),
    .C1(_05336_),
    .X(_05337_));
 sky130_fd_sc_hd__a22o_2 _08162_ (.A1(\tag_array.dirty0[5] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\tag_array.dirty0[6] ),
    .X(_05338_));
 sky130_fd_sc_hd__a221o_2 _08163_ (.A1(\tag_array.dirty0[4] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\tag_array.dirty0[7] ),
    .C1(_05338_),
    .X(_05339_));
 sky130_fd_sc_hd__a22o_2 _08164_ (.A1(_03522_),
    .A2(_05333_),
    .B1(_05337_),
    .B2(_03506_),
    .X(_05340_));
 sky130_fd_sc_hd__a22o_2 _08165_ (.A1(_03518_),
    .A2(_05335_),
    .B1(_05339_),
    .B2(_03526_),
    .X(_05341_));
 sky130_fd_sc_hd__or2_2 _08166_ (.A(_05340_),
    .B(_05341_),
    .X(_00129_));
 sky130_fd_sc_hd__a22o_2 _08167_ (.A1(\lru_array.lru_mem[13] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\lru_array.lru_mem[14] ),
    .X(_05342_));
 sky130_fd_sc_hd__a221o_2 _08168_ (.A1(\lru_array.lru_mem[12] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\lru_array.lru_mem[15] ),
    .C1(_05342_),
    .X(_05343_));
 sky130_fd_sc_hd__a22o_2 _08169_ (.A1(\lru_array.lru_mem[5] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\lru_array.lru_mem[6] ),
    .X(_05344_));
 sky130_fd_sc_hd__a221o_2 _08170_ (.A1(\lru_array.lru_mem[4] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\lru_array.lru_mem[7] ),
    .C1(_05344_),
    .X(_05345_));
 sky130_fd_sc_hd__a22o_2 _08171_ (.A1(\lru_array.lru_mem[9] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\lru_array.lru_mem[10] ),
    .X(_05346_));
 sky130_fd_sc_hd__a221o_2 _08172_ (.A1(\lru_array.lru_mem[8] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\lru_array.lru_mem[11] ),
    .C1(_05346_),
    .X(_05347_));
 sky130_fd_sc_hd__a22o_2 _08173_ (.A1(\lru_array.lru_mem[1] ),
    .A2(_03508_),
    .B1(_03510_),
    .B2(\lru_array.lru_mem[2] ),
    .X(_05348_));
 sky130_fd_sc_hd__a221o_2 _08174_ (.A1(\lru_array.lru_mem[0] ),
    .A2(_03513_),
    .B1(_03515_),
    .B2(\lru_array.lru_mem[3] ),
    .C1(_05348_),
    .X(_05349_));
 sky130_fd_sc_hd__a22o_2 _08175_ (.A1(_03522_),
    .A2(_05343_),
    .B1(_05347_),
    .B2(_03506_),
    .X(_05350_));
 sky130_fd_sc_hd__a22o_2 _08176_ (.A1(_03526_),
    .A2(_05345_),
    .B1(_05349_),
    .B2(_03518_),
    .X(_05351_));
 sky130_fd_sc_hd__or2_2 _08177_ (.A(_05350_),
    .B(_05351_),
    .X(_00128_));
 sky130_fd_sc_hd__and3_2 _08178_ (.A(\fsm.state[3] ),
    .B(_03213_),
    .C(_03285_),
    .X(_00185_));
 sky130_fd_sc_hd__a21boi_2 _08179_ (.A1(_03213_),
    .A2(_03285_),
    .B1_N(\fsm.state[3] ),
    .Y(_00183_));
 sky130_fd_sc_hd__o21a_2 _08180_ (.A1(cpu_write),
    .A2(cpu_read),
    .B1(\fsm.state[0] ),
    .X(_00184_));
 sky130_fd_sc_hd__nor2_2 _08181_ (.A(_03511_),
    .B(_03519_),
    .Y(_05352_));
 sky130_fd_sc_hd__o31ai_2 _08182_ (.A1(_03146_),
    .A2(_03333_),
    .A3(_03347_),
    .B1(cpu_ready),
    .Y(_05353_));
 sky130_fd_sc_hd__or3_2 _08183_ (.A(_03511_),
    .B(_03519_),
    .C(_05353_),
    .X(_05354_));
 sky130_fd_sc_hd__nor2_2 _08184_ (.A(\fsm.lru_out ),
    .B(_03147_),
    .Y(_05355_));
 sky130_fd_sc_hd__a21o_2 _08185_ (.A1(\fsm.state[2] ),
    .A2(_03236_),
    .B1(_05355_),
    .X(_05356_));
 sky130_fd_sc_hd__mux2_1 _08186_ (.A0(_05356_),
    .A1(\lru_array.lru_mem[2] ),
    .S(_05354_),
    .X(_00195_));
 sky130_fd_sc_hd__and3_2 _08187_ (.A(mem_ready),
    .B(mem_read),
    .C(\fsm.lru_out ),
    .X(_05357_));
 sky130_fd_sc_hd__o41a_2 _08188_ (.A1(_03320_),
    .A2(_03326_),
    .A3(_03327_),
    .A4(_03332_),
    .B1(\fsm.state[2] ),
    .X(_05358_));
 sky130_fd_sc_hd__and3_2 _08189_ (.A(cpu_write),
    .B(_03315_),
    .C(_05358_),
    .X(_05359_));
 sky130_fd_sc_hd__a31o_2 _08190_ (.A1(cpu_write),
    .A2(_03347_),
    .A3(_05358_),
    .B1(_05357_),
    .X(_05360_));
 sky130_fd_sc_hd__nand2_2 _08191_ (.A(_03515_),
    .B(_03526_),
    .Y(_05361_));
 sky130_fd_sc_hd__nand2b_2 _08192_ (.A_N(_05361_),
    .B(_05360_),
    .Y(_05362_));
 sky130_fd_sc_hd__and3_2 _08193_ (.A(mem_ready),
    .B(mem_read),
    .C(cpu_addr[7]),
    .X(_05363_));
 sky130_fd_sc_hd__and3_2 _08194_ (.A(\fsm.state[2] ),
    .B(cpu_write),
    .C(_03236_),
    .X(_05364_));
 sky130_fd_sc_hd__a221o_2 _08195_ (.A1(\fsm.tag_out1[0] ),
    .A2(_05359_),
    .B1(_05364_),
    .B2(\fsm.tag_out0[0] ),
    .C1(_05363_),
    .X(_05365_));
 sky130_fd_sc_hd__mux2_1 _08196_ (.A0(_05365_),
    .A1(\tag_array.tag1[7][0] ),
    .S(_05362_),
    .X(_00196_));
 sky130_fd_sc_hd__nor2_2 _08197_ (.A(_03135_),
    .B(_03147_),
    .Y(_05366_));
 sky130_fd_sc_hd__a221o_2 _08198_ (.A1(\fsm.tag_out1[1] ),
    .A2(_05359_),
    .B1(_05364_),
    .B2(\fsm.tag_out0[1] ),
    .C1(_05366_),
    .X(_05367_));
 sky130_fd_sc_hd__mux2_1 _08199_ (.A0(_05367_),
    .A1(\tag_array.tag1[7][1] ),
    .S(_05362_),
    .X(_00197_));
 sky130_fd_sc_hd__nor2_2 _08200_ (.A(_03136_),
    .B(_03147_),
    .Y(_05368_));
 sky130_fd_sc_hd__a221o_2 _08201_ (.A1(\fsm.tag_out1[2] ),
    .A2(_05359_),
    .B1(_05364_),
    .B2(\fsm.tag_out0[2] ),
    .C1(_05368_),
    .X(_05369_));
 sky130_fd_sc_hd__mux2_1 _08202_ (.A0(_05369_),
    .A1(\tag_array.tag1[7][2] ),
    .S(_05362_),
    .X(_00198_));
 sky130_fd_sc_hd__and3_2 _08203_ (.A(mem_ready),
    .B(mem_read),
    .C(cpu_addr[10]),
    .X(_05370_));
 sky130_fd_sc_hd__a221o_2 _08204_ (.A1(\fsm.tag_out1[3] ),
    .A2(_05359_),
    .B1(_05364_),
    .B2(\fsm.tag_out0[3] ),
    .C1(_05370_),
    .X(_05371_));
 sky130_fd_sc_hd__mux2_1 _08205_ (.A0(_05371_),
    .A1(\tag_array.tag1[7][3] ),
    .S(_05362_),
    .X(_00199_));
 sky130_fd_sc_hd__and3_2 _08206_ (.A(mem_ready),
    .B(mem_read),
    .C(cpu_addr[11]),
    .X(_05372_));
 sky130_fd_sc_hd__a221o_2 _08207_ (.A1(\fsm.tag_out1[4] ),
    .A2(_05359_),
    .B1(_05364_),
    .B2(\fsm.tag_out0[4] ),
    .C1(_05372_),
    .X(_05373_));
 sky130_fd_sc_hd__mux2_1 _08208_ (.A0(_05373_),
    .A1(\tag_array.tag1[7][4] ),
    .S(_05362_),
    .X(_00200_));
 sky130_fd_sc_hd__and3_2 _08209_ (.A(mem_ready),
    .B(mem_read),
    .C(cpu_addr[12]),
    .X(_05374_));
 sky130_fd_sc_hd__a221o_2 _08210_ (.A1(\fsm.tag_out1[5] ),
    .A2(_05359_),
    .B1(_05364_),
    .B2(\fsm.tag_out0[5] ),
    .C1(_05374_),
    .X(_05375_));
 sky130_fd_sc_hd__mux2_1 _08211_ (.A0(_05375_),
    .A1(\tag_array.tag1[7][5] ),
    .S(_05362_),
    .X(_00201_));
 sky130_fd_sc_hd__and3_2 _08212_ (.A(mem_ready),
    .B(mem_read),
    .C(cpu_addr[13]),
    .X(_05376_));
 sky130_fd_sc_hd__a221o_2 _08213_ (.A1(\fsm.tag_out1[6] ),
    .A2(_05359_),
    .B1(_05364_),
    .B2(\fsm.tag_out0[6] ),
    .C1(_05376_),
    .X(_05377_));
 sky130_fd_sc_hd__mux2_1 _08214_ (.A0(_05377_),
    .A1(\tag_array.tag1[7][6] ),
    .S(_05362_),
    .X(_00202_));
 sky130_fd_sc_hd__and3_2 _08215_ (.A(mem_ready),
    .B(mem_read),
    .C(cpu_addr[14]),
    .X(_05378_));
 sky130_fd_sc_hd__a221o_2 _08216_ (.A1(\fsm.tag_out1[7] ),
    .A2(_05359_),
    .B1(_05364_),
    .B2(\fsm.tag_out0[7] ),
    .C1(_05378_),
    .X(_05379_));
 sky130_fd_sc_hd__mux2_1 _08217_ (.A0(_05379_),
    .A1(\tag_array.tag1[7][7] ),
    .S(_05362_),
    .X(_00203_));
 sky130_fd_sc_hd__and3_2 _08218_ (.A(mem_ready),
    .B(mem_read),
    .C(cpu_addr[15]),
    .X(_05380_));
 sky130_fd_sc_hd__a221o_2 _08219_ (.A1(\fsm.tag_out1[8] ),
    .A2(_05359_),
    .B1(_05364_),
    .B2(\fsm.tag_out0[8] ),
    .C1(_05380_),
    .X(_05381_));
 sky130_fd_sc_hd__mux2_1 _08220_ (.A0(_05381_),
    .A1(\tag_array.tag1[7][8] ),
    .S(_05362_),
    .X(_00204_));
 sky130_fd_sc_hd__and3_2 _08221_ (.A(mem_ready),
    .B(mem_read),
    .C(cpu_addr[16]),
    .X(_05382_));
 sky130_fd_sc_hd__a221o_2 _08222_ (.A1(\fsm.tag_out1[9] ),
    .A2(_05359_),
    .B1(_05364_),
    .B2(\fsm.tag_out0[9] ),
    .C1(_05382_),
    .X(_05383_));
 sky130_fd_sc_hd__mux2_1 _08223_ (.A0(_05383_),
    .A1(\tag_array.tag1[7][9] ),
    .S(_05362_),
    .X(_00205_));
 sky130_fd_sc_hd__and3_2 _08224_ (.A(mem_ready),
    .B(mem_read),
    .C(cpu_addr[17]),
    .X(_05384_));
 sky130_fd_sc_hd__a221o_2 _08225_ (.A1(\fsm.tag_out1[10] ),
    .A2(_05359_),
    .B1(_05364_),
    .B2(\fsm.tag_out0[10] ),
    .C1(_05384_),
    .X(_05385_));
 sky130_fd_sc_hd__mux2_1 _08226_ (.A0(_05385_),
    .A1(\tag_array.tag1[7][10] ),
    .S(_05362_),
    .X(_00206_));
 sky130_fd_sc_hd__nor2_2 _08227_ (.A(_03139_),
    .B(_03147_),
    .Y(_05386_));
 sky130_fd_sc_hd__a221o_2 _08228_ (.A1(\fsm.tag_out1[11] ),
    .A2(_05359_),
    .B1(_05364_),
    .B2(\fsm.tag_out0[11] ),
    .C1(_05386_),
    .X(_05387_));
 sky130_fd_sc_hd__mux2_1 _08229_ (.A0(_05387_),
    .A1(\tag_array.tag1[7][11] ),
    .S(_05362_),
    .X(_00207_));
 sky130_fd_sc_hd__and3_2 _08230_ (.A(mem_ready),
    .B(mem_read),
    .C(cpu_addr[19]),
    .X(_05388_));
 sky130_fd_sc_hd__a221o_2 _08231_ (.A1(\fsm.tag_out1[12] ),
    .A2(_05359_),
    .B1(_05364_),
    .B2(\fsm.tag_out0[12] ),
    .C1(_05388_),
    .X(_05389_));
 sky130_fd_sc_hd__mux2_1 _08232_ (.A0(_05389_),
    .A1(\tag_array.tag1[7][12] ),
    .S(_05362_),
    .X(_00208_));
 sky130_fd_sc_hd__and3_2 _08233_ (.A(mem_ready),
    .B(mem_read),
    .C(cpu_addr[20]),
    .X(_05390_));
 sky130_fd_sc_hd__a221o_2 _08234_ (.A1(\fsm.tag_out1[13] ),
    .A2(_05359_),
    .B1(_05364_),
    .B2(\fsm.tag_out0[13] ),
    .C1(_05390_),
    .X(_05391_));
 sky130_fd_sc_hd__mux2_1 _08235_ (.A0(_05391_),
    .A1(\tag_array.tag1[7][13] ),
    .S(_05362_),
    .X(_00209_));
 sky130_fd_sc_hd__nor2_2 _08236_ (.A(_03140_),
    .B(_03147_),
    .Y(_05392_));
 sky130_fd_sc_hd__a221o_2 _08237_ (.A1(\fsm.tag_out1[14] ),
    .A2(_05359_),
    .B1(_05364_),
    .B2(\fsm.tag_out0[14] ),
    .C1(_05392_),
    .X(_05393_));
 sky130_fd_sc_hd__mux2_1 _08238_ (.A0(_05393_),
    .A1(\tag_array.tag1[7][14] ),
    .S(_05362_),
    .X(_00210_));
 sky130_fd_sc_hd__and3_2 _08239_ (.A(mem_ready),
    .B(mem_read),
    .C(cpu_addr[22]),
    .X(_05394_));
 sky130_fd_sc_hd__a221o_2 _08240_ (.A1(\fsm.tag_out1[15] ),
    .A2(_05359_),
    .B1(_05364_),
    .B2(\fsm.tag_out0[15] ),
    .C1(_05394_),
    .X(_05395_));
 sky130_fd_sc_hd__mux2_1 _08241_ (.A0(_05395_),
    .A1(\tag_array.tag1[7][15] ),
    .S(_05362_),
    .X(_00211_));
 sky130_fd_sc_hd__and3_2 _08242_ (.A(mem_ready),
    .B(mem_read),
    .C(cpu_addr[23]),
    .X(_05396_));
 sky130_fd_sc_hd__a221o_2 _08243_ (.A1(\fsm.tag_out1[16] ),
    .A2(_05359_),
    .B1(_05364_),
    .B2(\fsm.tag_out0[16] ),
    .C1(_05396_),
    .X(_05397_));
 sky130_fd_sc_hd__mux2_1 _08244_ (.A0(_05397_),
    .A1(\tag_array.tag1[7][16] ),
    .S(_05362_),
    .X(_00212_));
 sky130_fd_sc_hd__and3_2 _08245_ (.A(mem_ready),
    .B(mem_read),
    .C(cpu_addr[24]),
    .X(_05398_));
 sky130_fd_sc_hd__a221o_2 _08246_ (.A1(\fsm.tag_out1[17] ),
    .A2(_05359_),
    .B1(_05364_),
    .B2(\fsm.tag_out0[17] ),
    .C1(_05398_),
    .X(_05399_));
 sky130_fd_sc_hd__mux2_1 _08247_ (.A0(_05399_),
    .A1(\tag_array.tag1[7][17] ),
    .S(_05362_),
    .X(_00213_));
 sky130_fd_sc_hd__nor2_2 _08248_ (.A(_03142_),
    .B(_03147_),
    .Y(_05400_));
 sky130_fd_sc_hd__a221o_2 _08249_ (.A1(\fsm.tag_out1[18] ),
    .A2(_05359_),
    .B1(_05364_),
    .B2(\fsm.tag_out0[18] ),
    .C1(_05400_),
    .X(_05401_));
 sky130_fd_sc_hd__mux2_1 _08250_ (.A0(_05401_),
    .A1(\tag_array.tag1[7][18] ),
    .S(_05362_),
    .X(_00214_));
 sky130_fd_sc_hd__and3_2 _08251_ (.A(mem_ready),
    .B(mem_read),
    .C(cpu_addr[26]),
    .X(_05402_));
 sky130_fd_sc_hd__a221o_2 _08252_ (.A1(\fsm.tag_out1[19] ),
    .A2(_05359_),
    .B1(_05364_),
    .B2(\fsm.tag_out0[19] ),
    .C1(_05402_),
    .X(_05403_));
 sky130_fd_sc_hd__mux2_1 _08253_ (.A0(_05403_),
    .A1(\tag_array.tag1[7][19] ),
    .S(_05362_),
    .X(_00215_));
 sky130_fd_sc_hd__nor2_2 _08254_ (.A(_03143_),
    .B(_03147_),
    .Y(_05404_));
 sky130_fd_sc_hd__a221o_2 _08255_ (.A1(\fsm.tag_out1[20] ),
    .A2(_05359_),
    .B1(_05364_),
    .B2(\fsm.tag_out0[20] ),
    .C1(_05404_),
    .X(_05405_));
 sky130_fd_sc_hd__mux2_1 _08256_ (.A0(_05405_),
    .A1(\tag_array.tag1[7][20] ),
    .S(_05362_),
    .X(_00216_));
 sky130_fd_sc_hd__and3_2 _08257_ (.A(mem_ready),
    .B(mem_read),
    .C(cpu_addr[28]),
    .X(_05406_));
 sky130_fd_sc_hd__a221o_2 _08258_ (.A1(\fsm.tag_out1[21] ),
    .A2(_05359_),
    .B1(_05364_),
    .B2(\fsm.tag_out0[21] ),
    .C1(_05406_),
    .X(_05407_));
 sky130_fd_sc_hd__mux2_1 _08259_ (.A0(_05407_),
    .A1(\tag_array.tag1[7][21] ),
    .S(_05362_),
    .X(_00217_));
 sky130_fd_sc_hd__and3_2 _08260_ (.A(mem_ready),
    .B(mem_read),
    .C(cpu_addr[29]),
    .X(_05408_));
 sky130_fd_sc_hd__a221o_2 _08261_ (.A1(\fsm.tag_out1[22] ),
    .A2(_05359_),
    .B1(_05364_),
    .B2(\fsm.tag_out0[22] ),
    .C1(_05408_),
    .X(_05409_));
 sky130_fd_sc_hd__mux2_1 _08262_ (.A0(_05409_),
    .A1(\tag_array.tag1[7][22] ),
    .S(_05362_),
    .X(_00218_));
 sky130_fd_sc_hd__and3_2 _08263_ (.A(mem_ready),
    .B(mem_read),
    .C(cpu_addr[30]),
    .X(_05410_));
 sky130_fd_sc_hd__a221o_2 _08264_ (.A1(\fsm.tag_out1[23] ),
    .A2(_05359_),
    .B1(_05364_),
    .B2(\fsm.tag_out0[23] ),
    .C1(_05410_),
    .X(_05411_));
 sky130_fd_sc_hd__mux2_1 _08265_ (.A0(_05411_),
    .A1(\tag_array.tag1[7][23] ),
    .S(_05362_),
    .X(_00219_));
 sky130_fd_sc_hd__and3_2 _08266_ (.A(mem_ready),
    .B(mem_read),
    .C(cpu_addr[31]),
    .X(_05412_));
 sky130_fd_sc_hd__a221o_2 _08267_ (.A1(\fsm.tag_out1[24] ),
    .A2(_05359_),
    .B1(_05364_),
    .B2(\fsm.tag_out0[24] ),
    .C1(_05412_),
    .X(_05413_));
 sky130_fd_sc_hd__mux2_1 _08268_ (.A0(_05413_),
    .A1(\tag_array.tag1[7][24] ),
    .S(_05362_),
    .X(_00220_));
 sky130_fd_sc_hd__a31oi_2 _08269_ (.A1(\fsm.state[2] ),
    .A2(cpu_write),
    .A3(_03236_),
    .B1(_05355_),
    .Y(_05414_));
 sky130_fd_sc_hd__a31o_2 _08270_ (.A1(\fsm.state[2] ),
    .A2(cpu_write),
    .A3(_03236_),
    .B1(_05355_),
    .X(_05415_));
 sky130_fd_sc_hd__nor2_2 _08271_ (.A(_03514_),
    .B(_03519_),
    .Y(_05416_));
 sky130_fd_sc_hd__and2_2 _08272_ (.A(_05415_),
    .B(_05416_),
    .X(_05417_));
 sky130_fd_sc_hd__or2_2 _08273_ (.A(mem_read),
    .B(\fsm.state[2] ),
    .X(_05418_));
 sky130_fd_sc_hd__mux2_1 _08274_ (.A0(mem_rdata[0]),
    .A1(cpu_wdata[0]),
    .S(cpu_write),
    .X(_05419_));
 sky130_fd_sc_hd__and2_2 _08275_ (.A(_05418_),
    .B(_05419_),
    .X(_05420_));
 sky130_fd_sc_hd__mux2_1 _08276_ (.A0(\data_array.data0[0][0] ),
    .A1(_05420_),
    .S(_05417_),
    .X(_00221_));
 sky130_fd_sc_hd__mux2_1 _08277_ (.A0(mem_rdata[1]),
    .A1(cpu_wdata[1]),
    .S(cpu_write),
    .X(_05421_));
 sky130_fd_sc_hd__and2_2 _08278_ (.A(_05418_),
    .B(_05421_),
    .X(_05422_));
 sky130_fd_sc_hd__mux2_1 _08279_ (.A0(\data_array.data0[0][1] ),
    .A1(_05422_),
    .S(_05417_),
    .X(_00222_));
 sky130_fd_sc_hd__mux2_1 _08280_ (.A0(mem_rdata[2]),
    .A1(cpu_wdata[2]),
    .S(cpu_write),
    .X(_05423_));
 sky130_fd_sc_hd__and2_2 _08281_ (.A(_05418_),
    .B(_05423_),
    .X(_05424_));
 sky130_fd_sc_hd__mux2_1 _08282_ (.A0(\data_array.data0[0][2] ),
    .A1(_05424_),
    .S(_05417_),
    .X(_00223_));
 sky130_fd_sc_hd__mux2_1 _08283_ (.A0(mem_rdata[3]),
    .A1(cpu_wdata[3]),
    .S(cpu_write),
    .X(_05425_));
 sky130_fd_sc_hd__and2_2 _08284_ (.A(_05418_),
    .B(_05425_),
    .X(_05426_));
 sky130_fd_sc_hd__mux2_1 _08285_ (.A0(\data_array.data0[0][3] ),
    .A1(_05426_),
    .S(_05417_),
    .X(_00224_));
 sky130_fd_sc_hd__mux2_1 _08286_ (.A0(mem_rdata[4]),
    .A1(cpu_wdata[4]),
    .S(cpu_write),
    .X(_05427_));
 sky130_fd_sc_hd__and2_2 _08287_ (.A(_05418_),
    .B(_05427_),
    .X(_05428_));
 sky130_fd_sc_hd__mux2_1 _08288_ (.A0(\data_array.data0[0][4] ),
    .A1(_05428_),
    .S(_05417_),
    .X(_00225_));
 sky130_fd_sc_hd__mux2_1 _08289_ (.A0(mem_rdata[5]),
    .A1(cpu_wdata[5]),
    .S(cpu_write),
    .X(_05429_));
 sky130_fd_sc_hd__and2_2 _08290_ (.A(_05418_),
    .B(_05429_),
    .X(_05430_));
 sky130_fd_sc_hd__mux2_1 _08291_ (.A0(\data_array.data0[0][5] ),
    .A1(_05430_),
    .S(_05417_),
    .X(_00226_));
 sky130_fd_sc_hd__mux2_1 _08292_ (.A0(mem_rdata[6]),
    .A1(cpu_wdata[6]),
    .S(cpu_write),
    .X(_05431_));
 sky130_fd_sc_hd__and2_2 _08293_ (.A(_05418_),
    .B(_05431_),
    .X(_05432_));
 sky130_fd_sc_hd__mux2_1 _08294_ (.A0(\data_array.data0[0][6] ),
    .A1(_05432_),
    .S(_05417_),
    .X(_00227_));
 sky130_fd_sc_hd__mux2_1 _08295_ (.A0(mem_rdata[7]),
    .A1(cpu_wdata[7]),
    .S(cpu_write),
    .X(_05433_));
 sky130_fd_sc_hd__and2_2 _08296_ (.A(_05418_),
    .B(_05433_),
    .X(_05434_));
 sky130_fd_sc_hd__mux2_1 _08297_ (.A0(\data_array.data0[0][7] ),
    .A1(_05434_),
    .S(_05417_),
    .X(_00228_));
 sky130_fd_sc_hd__mux2_1 _08298_ (.A0(mem_rdata[8]),
    .A1(cpu_wdata[8]),
    .S(cpu_write),
    .X(_05435_));
 sky130_fd_sc_hd__and2_2 _08299_ (.A(_05418_),
    .B(_05435_),
    .X(_05436_));
 sky130_fd_sc_hd__mux2_1 _08300_ (.A0(\data_array.data0[0][8] ),
    .A1(_05436_),
    .S(_05417_),
    .X(_00229_));
 sky130_fd_sc_hd__mux2_1 _08301_ (.A0(mem_rdata[9]),
    .A1(cpu_wdata[9]),
    .S(cpu_write),
    .X(_05437_));
 sky130_fd_sc_hd__and2_2 _08302_ (.A(_05418_),
    .B(_05437_),
    .X(_05438_));
 sky130_fd_sc_hd__mux2_1 _08303_ (.A0(\data_array.data0[0][9] ),
    .A1(_05438_),
    .S(_05417_),
    .X(_00230_));
 sky130_fd_sc_hd__mux2_1 _08304_ (.A0(mem_rdata[10]),
    .A1(cpu_wdata[10]),
    .S(cpu_write),
    .X(_05439_));
 sky130_fd_sc_hd__and2_2 _08305_ (.A(_05418_),
    .B(_05439_),
    .X(_05440_));
 sky130_fd_sc_hd__mux2_1 _08306_ (.A0(\data_array.data0[0][10] ),
    .A1(_05440_),
    .S(_05417_),
    .X(_00231_));
 sky130_fd_sc_hd__mux2_1 _08307_ (.A0(mem_rdata[11]),
    .A1(cpu_wdata[11]),
    .S(cpu_write),
    .X(_05441_));
 sky130_fd_sc_hd__and2_2 _08308_ (.A(_05418_),
    .B(_05441_),
    .X(_05442_));
 sky130_fd_sc_hd__mux2_1 _08309_ (.A0(\data_array.data0[0][11] ),
    .A1(_05442_),
    .S(_05417_),
    .X(_00232_));
 sky130_fd_sc_hd__mux2_1 _08310_ (.A0(mem_rdata[12]),
    .A1(cpu_wdata[12]),
    .S(cpu_write),
    .X(_05443_));
 sky130_fd_sc_hd__and2_2 _08311_ (.A(_05418_),
    .B(_05443_),
    .X(_05444_));
 sky130_fd_sc_hd__mux2_1 _08312_ (.A0(\data_array.data0[0][12] ),
    .A1(_05444_),
    .S(_05417_),
    .X(_00233_));
 sky130_fd_sc_hd__mux2_1 _08313_ (.A0(mem_rdata[13]),
    .A1(cpu_wdata[13]),
    .S(cpu_write),
    .X(_05445_));
 sky130_fd_sc_hd__and2_2 _08314_ (.A(_05418_),
    .B(_05445_),
    .X(_05446_));
 sky130_fd_sc_hd__mux2_1 _08315_ (.A0(\data_array.data0[0][13] ),
    .A1(_05446_),
    .S(_05417_),
    .X(_00234_));
 sky130_fd_sc_hd__mux2_1 _08316_ (.A0(mem_rdata[14]),
    .A1(cpu_wdata[14]),
    .S(cpu_write),
    .X(_05447_));
 sky130_fd_sc_hd__and2_2 _08317_ (.A(_05418_),
    .B(_05447_),
    .X(_05448_));
 sky130_fd_sc_hd__mux2_1 _08318_ (.A0(\data_array.data0[0][14] ),
    .A1(_05448_),
    .S(_05417_),
    .X(_00235_));
 sky130_fd_sc_hd__mux2_1 _08319_ (.A0(mem_rdata[15]),
    .A1(cpu_wdata[15]),
    .S(cpu_write),
    .X(_05449_));
 sky130_fd_sc_hd__and2_2 _08320_ (.A(_05418_),
    .B(_05449_),
    .X(_05450_));
 sky130_fd_sc_hd__mux2_1 _08321_ (.A0(\data_array.data0[0][15] ),
    .A1(_05450_),
    .S(_05417_),
    .X(_00236_));
 sky130_fd_sc_hd__mux2_1 _08322_ (.A0(mem_rdata[16]),
    .A1(cpu_wdata[16]),
    .S(cpu_write),
    .X(_05451_));
 sky130_fd_sc_hd__and2_2 _08323_ (.A(_05418_),
    .B(_05451_),
    .X(_05452_));
 sky130_fd_sc_hd__mux2_1 _08324_ (.A0(\data_array.data0[0][16] ),
    .A1(_05452_),
    .S(_05417_),
    .X(_00237_));
 sky130_fd_sc_hd__mux2_1 _08325_ (.A0(mem_rdata[17]),
    .A1(cpu_wdata[17]),
    .S(cpu_write),
    .X(_05453_));
 sky130_fd_sc_hd__and2_2 _08326_ (.A(_05418_),
    .B(_05453_),
    .X(_05454_));
 sky130_fd_sc_hd__mux2_1 _08327_ (.A0(\data_array.data0[0][17] ),
    .A1(_05454_),
    .S(_05417_),
    .X(_00238_));
 sky130_fd_sc_hd__mux2_1 _08328_ (.A0(mem_rdata[18]),
    .A1(cpu_wdata[18]),
    .S(cpu_write),
    .X(_05455_));
 sky130_fd_sc_hd__and2_2 _08329_ (.A(_05418_),
    .B(_05455_),
    .X(_05456_));
 sky130_fd_sc_hd__mux2_1 _08330_ (.A0(\data_array.data0[0][18] ),
    .A1(_05456_),
    .S(_05417_),
    .X(_00239_));
 sky130_fd_sc_hd__mux2_1 _08331_ (.A0(mem_rdata[19]),
    .A1(cpu_wdata[19]),
    .S(cpu_write),
    .X(_05457_));
 sky130_fd_sc_hd__and2_2 _08332_ (.A(_05418_),
    .B(_05457_),
    .X(_05458_));
 sky130_fd_sc_hd__mux2_1 _08333_ (.A0(\data_array.data0[0][19] ),
    .A1(_05458_),
    .S(_05417_),
    .X(_00240_));
 sky130_fd_sc_hd__mux2_1 _08334_ (.A0(mem_rdata[20]),
    .A1(cpu_wdata[20]),
    .S(cpu_write),
    .X(_05459_));
 sky130_fd_sc_hd__and2_2 _08335_ (.A(_05418_),
    .B(_05459_),
    .X(_05460_));
 sky130_fd_sc_hd__mux2_1 _08336_ (.A0(\data_array.data0[0][20] ),
    .A1(_05460_),
    .S(_05417_),
    .X(_00241_));
 sky130_fd_sc_hd__mux2_1 _08337_ (.A0(mem_rdata[21]),
    .A1(cpu_wdata[21]),
    .S(cpu_write),
    .X(_05461_));
 sky130_fd_sc_hd__and2_2 _08338_ (.A(_05418_),
    .B(_05461_),
    .X(_05462_));
 sky130_fd_sc_hd__mux2_1 _08339_ (.A0(\data_array.data0[0][21] ),
    .A1(_05462_),
    .S(_05417_),
    .X(_00242_));
 sky130_fd_sc_hd__mux2_1 _08340_ (.A0(mem_rdata[22]),
    .A1(cpu_wdata[22]),
    .S(cpu_write),
    .X(_05463_));
 sky130_fd_sc_hd__and2_2 _08341_ (.A(_05418_),
    .B(_05463_),
    .X(_05464_));
 sky130_fd_sc_hd__mux2_1 _08342_ (.A0(\data_array.data0[0][22] ),
    .A1(_05464_),
    .S(_05417_),
    .X(_00243_));
 sky130_fd_sc_hd__mux2_1 _08343_ (.A0(mem_rdata[23]),
    .A1(cpu_wdata[23]),
    .S(cpu_write),
    .X(_05465_));
 sky130_fd_sc_hd__and2_2 _08344_ (.A(_05418_),
    .B(_05465_),
    .X(_05466_));
 sky130_fd_sc_hd__mux2_1 _08345_ (.A0(\data_array.data0[0][23] ),
    .A1(_05466_),
    .S(_05417_),
    .X(_00244_));
 sky130_fd_sc_hd__mux2_1 _08346_ (.A0(mem_rdata[24]),
    .A1(cpu_wdata[24]),
    .S(cpu_write),
    .X(_05467_));
 sky130_fd_sc_hd__and2_2 _08347_ (.A(_05418_),
    .B(_05467_),
    .X(_05468_));
 sky130_fd_sc_hd__mux2_1 _08348_ (.A0(\data_array.data0[0][24] ),
    .A1(_05468_),
    .S(_05417_),
    .X(_00245_));
 sky130_fd_sc_hd__mux2_1 _08349_ (.A0(mem_rdata[25]),
    .A1(cpu_wdata[25]),
    .S(cpu_write),
    .X(_05469_));
 sky130_fd_sc_hd__and2_2 _08350_ (.A(_05418_),
    .B(_05469_),
    .X(_05470_));
 sky130_fd_sc_hd__mux2_1 _08351_ (.A0(\data_array.data0[0][25] ),
    .A1(_05470_),
    .S(_05417_),
    .X(_00246_));
 sky130_fd_sc_hd__mux2_1 _08352_ (.A0(mem_rdata[26]),
    .A1(cpu_wdata[26]),
    .S(cpu_write),
    .X(_05471_));
 sky130_fd_sc_hd__and2_2 _08353_ (.A(_05418_),
    .B(_05471_),
    .X(_05472_));
 sky130_fd_sc_hd__mux2_1 _08354_ (.A0(\data_array.data0[0][26] ),
    .A1(_05472_),
    .S(_05417_),
    .X(_00247_));
 sky130_fd_sc_hd__mux2_1 _08355_ (.A0(mem_rdata[27]),
    .A1(cpu_wdata[27]),
    .S(cpu_write),
    .X(_05473_));
 sky130_fd_sc_hd__and2_2 _08356_ (.A(_05418_),
    .B(_05473_),
    .X(_05474_));
 sky130_fd_sc_hd__mux2_1 _08357_ (.A0(\data_array.data0[0][27] ),
    .A1(_05474_),
    .S(_05417_),
    .X(_00248_));
 sky130_fd_sc_hd__mux2_1 _08358_ (.A0(mem_rdata[28]),
    .A1(cpu_wdata[28]),
    .S(cpu_write),
    .X(_05475_));
 sky130_fd_sc_hd__and2_2 _08359_ (.A(_05418_),
    .B(_05475_),
    .X(_05476_));
 sky130_fd_sc_hd__mux2_1 _08360_ (.A0(\data_array.data0[0][28] ),
    .A1(_05476_),
    .S(_05417_),
    .X(_00249_));
 sky130_fd_sc_hd__mux2_1 _08361_ (.A0(mem_rdata[29]),
    .A1(cpu_wdata[29]),
    .S(cpu_write),
    .X(_05477_));
 sky130_fd_sc_hd__and2_2 _08362_ (.A(_05418_),
    .B(_05477_),
    .X(_05478_));
 sky130_fd_sc_hd__mux2_1 _08363_ (.A0(\data_array.data0[0][29] ),
    .A1(_05478_),
    .S(_05417_),
    .X(_00250_));
 sky130_fd_sc_hd__mux2_1 _08364_ (.A0(mem_rdata[30]),
    .A1(cpu_wdata[30]),
    .S(cpu_write),
    .X(_05479_));
 sky130_fd_sc_hd__and2_2 _08365_ (.A(_05418_),
    .B(_05479_),
    .X(_05480_));
 sky130_fd_sc_hd__mux2_1 _08366_ (.A0(\data_array.data0[0][30] ),
    .A1(_05480_),
    .S(_05417_),
    .X(_00251_));
 sky130_fd_sc_hd__mux2_1 _08367_ (.A0(mem_rdata[31]),
    .A1(cpu_wdata[31]),
    .S(cpu_write),
    .X(_05481_));
 sky130_fd_sc_hd__and2_2 _08368_ (.A(_05418_),
    .B(_05481_),
    .X(_05482_));
 sky130_fd_sc_hd__mux2_1 _08369_ (.A0(\data_array.data0[0][31] ),
    .A1(_05482_),
    .S(_05417_),
    .X(_00252_));
 sky130_fd_sc_hd__mux2_1 _08370_ (.A0(mem_rdata[32]),
    .A1(cpu_wdata[32]),
    .S(cpu_write),
    .X(_05483_));
 sky130_fd_sc_hd__and2_2 _08371_ (.A(_05418_),
    .B(_05483_),
    .X(_05484_));
 sky130_fd_sc_hd__mux2_1 _08372_ (.A0(\data_array.data0[0][32] ),
    .A1(_05484_),
    .S(_05417_),
    .X(_00253_));
 sky130_fd_sc_hd__mux2_1 _08373_ (.A0(mem_rdata[33]),
    .A1(cpu_wdata[33]),
    .S(cpu_write),
    .X(_05485_));
 sky130_fd_sc_hd__and2_2 _08374_ (.A(_05418_),
    .B(_05485_),
    .X(_05486_));
 sky130_fd_sc_hd__mux2_1 _08375_ (.A0(\data_array.data0[0][33] ),
    .A1(_05486_),
    .S(_05417_),
    .X(_00254_));
 sky130_fd_sc_hd__mux2_1 _08376_ (.A0(mem_rdata[34]),
    .A1(cpu_wdata[34]),
    .S(cpu_write),
    .X(_05487_));
 sky130_fd_sc_hd__and2_2 _08377_ (.A(_05418_),
    .B(_05487_),
    .X(_05488_));
 sky130_fd_sc_hd__mux2_1 _08378_ (.A0(\data_array.data0[0][34] ),
    .A1(_05488_),
    .S(_05417_),
    .X(_00255_));
 sky130_fd_sc_hd__mux2_1 _08379_ (.A0(mem_rdata[35]),
    .A1(cpu_wdata[35]),
    .S(cpu_write),
    .X(_05489_));
 sky130_fd_sc_hd__and2_2 _08380_ (.A(_05418_),
    .B(_05489_),
    .X(_05490_));
 sky130_fd_sc_hd__mux2_1 _08381_ (.A0(\data_array.data0[0][35] ),
    .A1(_05490_),
    .S(_05417_),
    .X(_00256_));
 sky130_fd_sc_hd__mux2_1 _08382_ (.A0(mem_rdata[36]),
    .A1(cpu_wdata[36]),
    .S(cpu_write),
    .X(_05491_));
 sky130_fd_sc_hd__and2_2 _08383_ (.A(_05418_),
    .B(_05491_),
    .X(_05492_));
 sky130_fd_sc_hd__mux2_1 _08384_ (.A0(\data_array.data0[0][36] ),
    .A1(_05492_),
    .S(_05417_),
    .X(_00257_));
 sky130_fd_sc_hd__mux2_1 _08385_ (.A0(mem_rdata[37]),
    .A1(cpu_wdata[37]),
    .S(cpu_write),
    .X(_05493_));
 sky130_fd_sc_hd__and2_2 _08386_ (.A(_05418_),
    .B(_05493_),
    .X(_05494_));
 sky130_fd_sc_hd__mux2_1 _08387_ (.A0(\data_array.data0[0][37] ),
    .A1(_05494_),
    .S(_05417_),
    .X(_00258_));
 sky130_fd_sc_hd__mux2_1 _08388_ (.A0(mem_rdata[38]),
    .A1(cpu_wdata[38]),
    .S(cpu_write),
    .X(_05495_));
 sky130_fd_sc_hd__and2_2 _08389_ (.A(_05418_),
    .B(_05495_),
    .X(_05496_));
 sky130_fd_sc_hd__mux2_1 _08390_ (.A0(\data_array.data0[0][38] ),
    .A1(_05496_),
    .S(_05417_),
    .X(_00259_));
 sky130_fd_sc_hd__mux2_1 _08391_ (.A0(mem_rdata[39]),
    .A1(cpu_wdata[39]),
    .S(cpu_write),
    .X(_05497_));
 sky130_fd_sc_hd__and2_2 _08392_ (.A(_05418_),
    .B(_05497_),
    .X(_05498_));
 sky130_fd_sc_hd__mux2_1 _08393_ (.A0(\data_array.data0[0][39] ),
    .A1(_05498_),
    .S(_05417_),
    .X(_00260_));
 sky130_fd_sc_hd__mux2_1 _08394_ (.A0(mem_rdata[40]),
    .A1(cpu_wdata[40]),
    .S(cpu_write),
    .X(_05499_));
 sky130_fd_sc_hd__and2_2 _08395_ (.A(_05418_),
    .B(_05499_),
    .X(_05500_));
 sky130_fd_sc_hd__mux2_1 _08396_ (.A0(\data_array.data0[0][40] ),
    .A1(_05500_),
    .S(_05417_),
    .X(_00261_));
 sky130_fd_sc_hd__mux2_1 _08397_ (.A0(mem_rdata[41]),
    .A1(cpu_wdata[41]),
    .S(cpu_write),
    .X(_05501_));
 sky130_fd_sc_hd__and2_2 _08398_ (.A(_05418_),
    .B(_05501_),
    .X(_05502_));
 sky130_fd_sc_hd__mux2_1 _08399_ (.A0(\data_array.data0[0][41] ),
    .A1(_05502_),
    .S(_05417_),
    .X(_00262_));
 sky130_fd_sc_hd__mux2_1 _08400_ (.A0(mem_rdata[42]),
    .A1(cpu_wdata[42]),
    .S(cpu_write),
    .X(_05503_));
 sky130_fd_sc_hd__and2_2 _08401_ (.A(_05418_),
    .B(_05503_),
    .X(_05504_));
 sky130_fd_sc_hd__mux2_1 _08402_ (.A0(\data_array.data0[0][42] ),
    .A1(_05504_),
    .S(_05417_),
    .X(_00263_));
 sky130_fd_sc_hd__mux2_1 _08403_ (.A0(mem_rdata[43]),
    .A1(cpu_wdata[43]),
    .S(cpu_write),
    .X(_05505_));
 sky130_fd_sc_hd__and2_2 _08404_ (.A(_05418_),
    .B(_05505_),
    .X(_05506_));
 sky130_fd_sc_hd__mux2_1 _08405_ (.A0(\data_array.data0[0][43] ),
    .A1(_05506_),
    .S(_05417_),
    .X(_00264_));
 sky130_fd_sc_hd__mux2_1 _08406_ (.A0(mem_rdata[44]),
    .A1(cpu_wdata[44]),
    .S(cpu_write),
    .X(_05507_));
 sky130_fd_sc_hd__and2_2 _08407_ (.A(_05418_),
    .B(_05507_),
    .X(_05508_));
 sky130_fd_sc_hd__mux2_1 _08408_ (.A0(\data_array.data0[0][44] ),
    .A1(_05508_),
    .S(_05417_),
    .X(_00265_));
 sky130_fd_sc_hd__mux2_1 _08409_ (.A0(mem_rdata[45]),
    .A1(cpu_wdata[45]),
    .S(cpu_write),
    .X(_05509_));
 sky130_fd_sc_hd__and2_2 _08410_ (.A(_05418_),
    .B(_05509_),
    .X(_05510_));
 sky130_fd_sc_hd__mux2_1 _08411_ (.A0(\data_array.data0[0][45] ),
    .A1(_05510_),
    .S(_05417_),
    .X(_00266_));
 sky130_fd_sc_hd__mux2_1 _08412_ (.A0(mem_rdata[46]),
    .A1(cpu_wdata[46]),
    .S(cpu_write),
    .X(_05511_));
 sky130_fd_sc_hd__and2_2 _08413_ (.A(_05418_),
    .B(_05511_),
    .X(_05512_));
 sky130_fd_sc_hd__mux2_1 _08414_ (.A0(\data_array.data0[0][46] ),
    .A1(_05512_),
    .S(_05417_),
    .X(_00267_));
 sky130_fd_sc_hd__mux2_1 _08415_ (.A0(mem_rdata[47]),
    .A1(cpu_wdata[47]),
    .S(cpu_write),
    .X(_05513_));
 sky130_fd_sc_hd__and2_2 _08416_ (.A(_05418_),
    .B(_05513_),
    .X(_05514_));
 sky130_fd_sc_hd__mux2_1 _08417_ (.A0(\data_array.data0[0][47] ),
    .A1(_05514_),
    .S(_05417_),
    .X(_00268_));
 sky130_fd_sc_hd__mux2_1 _08418_ (.A0(mem_rdata[48]),
    .A1(cpu_wdata[48]),
    .S(cpu_write),
    .X(_05515_));
 sky130_fd_sc_hd__and2_2 _08419_ (.A(_05418_),
    .B(_05515_),
    .X(_05516_));
 sky130_fd_sc_hd__mux2_1 _08420_ (.A0(\data_array.data0[0][48] ),
    .A1(_05516_),
    .S(_05417_),
    .X(_00269_));
 sky130_fd_sc_hd__mux2_1 _08421_ (.A0(mem_rdata[49]),
    .A1(cpu_wdata[49]),
    .S(cpu_write),
    .X(_05517_));
 sky130_fd_sc_hd__and2_2 _08422_ (.A(_05418_),
    .B(_05517_),
    .X(_05518_));
 sky130_fd_sc_hd__mux2_1 _08423_ (.A0(\data_array.data0[0][49] ),
    .A1(_05518_),
    .S(_05417_),
    .X(_00270_));
 sky130_fd_sc_hd__mux2_1 _08424_ (.A0(mem_rdata[50]),
    .A1(cpu_wdata[50]),
    .S(cpu_write),
    .X(_05519_));
 sky130_fd_sc_hd__and2_2 _08425_ (.A(_05418_),
    .B(_05519_),
    .X(_05520_));
 sky130_fd_sc_hd__mux2_1 _08426_ (.A0(\data_array.data0[0][50] ),
    .A1(_05520_),
    .S(_05417_),
    .X(_00271_));
 sky130_fd_sc_hd__mux2_1 _08427_ (.A0(mem_rdata[51]),
    .A1(cpu_wdata[51]),
    .S(cpu_write),
    .X(_05521_));
 sky130_fd_sc_hd__and2_2 _08428_ (.A(_05418_),
    .B(_05521_),
    .X(_05522_));
 sky130_fd_sc_hd__mux2_1 _08429_ (.A0(\data_array.data0[0][51] ),
    .A1(_05522_),
    .S(_05417_),
    .X(_00272_));
 sky130_fd_sc_hd__mux2_1 _08430_ (.A0(mem_rdata[52]),
    .A1(cpu_wdata[52]),
    .S(cpu_write),
    .X(_05523_));
 sky130_fd_sc_hd__and2_2 _08431_ (.A(_05418_),
    .B(_05523_),
    .X(_05524_));
 sky130_fd_sc_hd__mux2_1 _08432_ (.A0(\data_array.data0[0][52] ),
    .A1(_05524_),
    .S(_05417_),
    .X(_00273_));
 sky130_fd_sc_hd__mux2_1 _08433_ (.A0(mem_rdata[53]),
    .A1(cpu_wdata[53]),
    .S(cpu_write),
    .X(_05525_));
 sky130_fd_sc_hd__and2_2 _08434_ (.A(_05418_),
    .B(_05525_),
    .X(_05526_));
 sky130_fd_sc_hd__mux2_1 _08435_ (.A0(\data_array.data0[0][53] ),
    .A1(_05526_),
    .S(_05417_),
    .X(_00274_));
 sky130_fd_sc_hd__mux2_1 _08436_ (.A0(mem_rdata[54]),
    .A1(cpu_wdata[54]),
    .S(cpu_write),
    .X(_05527_));
 sky130_fd_sc_hd__and2_2 _08437_ (.A(_05418_),
    .B(_05527_),
    .X(_05528_));
 sky130_fd_sc_hd__mux2_1 _08438_ (.A0(\data_array.data0[0][54] ),
    .A1(_05528_),
    .S(_05417_),
    .X(_00275_));
 sky130_fd_sc_hd__mux2_1 _08439_ (.A0(mem_rdata[55]),
    .A1(cpu_wdata[55]),
    .S(cpu_write),
    .X(_05529_));
 sky130_fd_sc_hd__and2_2 _08440_ (.A(_05418_),
    .B(_05529_),
    .X(_05530_));
 sky130_fd_sc_hd__mux2_1 _08441_ (.A0(\data_array.data0[0][55] ),
    .A1(_05530_),
    .S(_05417_),
    .X(_00276_));
 sky130_fd_sc_hd__mux2_1 _08442_ (.A0(mem_rdata[56]),
    .A1(cpu_wdata[56]),
    .S(cpu_write),
    .X(_05531_));
 sky130_fd_sc_hd__and2_2 _08443_ (.A(_05418_),
    .B(_05531_),
    .X(_05532_));
 sky130_fd_sc_hd__mux2_1 _08444_ (.A0(\data_array.data0[0][56] ),
    .A1(_05532_),
    .S(_05417_),
    .X(_00277_));
 sky130_fd_sc_hd__mux2_1 _08445_ (.A0(mem_rdata[57]),
    .A1(cpu_wdata[57]),
    .S(cpu_write),
    .X(_05533_));
 sky130_fd_sc_hd__and2_2 _08446_ (.A(_05418_),
    .B(_05533_),
    .X(_05534_));
 sky130_fd_sc_hd__mux2_1 _08447_ (.A0(\data_array.data0[0][57] ),
    .A1(_05534_),
    .S(_05417_),
    .X(_00278_));
 sky130_fd_sc_hd__mux2_1 _08448_ (.A0(mem_rdata[58]),
    .A1(cpu_wdata[58]),
    .S(cpu_write),
    .X(_05535_));
 sky130_fd_sc_hd__and2_2 _08449_ (.A(_05418_),
    .B(_05535_),
    .X(_05536_));
 sky130_fd_sc_hd__mux2_1 _08450_ (.A0(\data_array.data0[0][58] ),
    .A1(_05536_),
    .S(_05417_),
    .X(_00279_));
 sky130_fd_sc_hd__mux2_1 _08451_ (.A0(mem_rdata[59]),
    .A1(cpu_wdata[59]),
    .S(cpu_write),
    .X(_05537_));
 sky130_fd_sc_hd__and2_2 _08452_ (.A(_05418_),
    .B(_05537_),
    .X(_05538_));
 sky130_fd_sc_hd__mux2_1 _08453_ (.A0(\data_array.data0[0][59] ),
    .A1(_05538_),
    .S(_05417_),
    .X(_00280_));
 sky130_fd_sc_hd__mux2_1 _08454_ (.A0(mem_rdata[60]),
    .A1(cpu_wdata[60]),
    .S(cpu_write),
    .X(_05539_));
 sky130_fd_sc_hd__and2_2 _08455_ (.A(_05418_),
    .B(_05539_),
    .X(_05540_));
 sky130_fd_sc_hd__mux2_1 _08456_ (.A0(\data_array.data0[0][60] ),
    .A1(_05540_),
    .S(_05417_),
    .X(_00281_));
 sky130_fd_sc_hd__mux2_1 _08457_ (.A0(mem_rdata[61]),
    .A1(cpu_wdata[61]),
    .S(cpu_write),
    .X(_05541_));
 sky130_fd_sc_hd__and2_2 _08458_ (.A(_05418_),
    .B(_05541_),
    .X(_05542_));
 sky130_fd_sc_hd__mux2_1 _08459_ (.A0(\data_array.data0[0][61] ),
    .A1(_05542_),
    .S(_05417_),
    .X(_00282_));
 sky130_fd_sc_hd__mux2_1 _08460_ (.A0(mem_rdata[62]),
    .A1(cpu_wdata[62]),
    .S(cpu_write),
    .X(_05543_));
 sky130_fd_sc_hd__and2_2 _08461_ (.A(_05418_),
    .B(_05543_),
    .X(_05544_));
 sky130_fd_sc_hd__mux2_1 _08462_ (.A0(\data_array.data0[0][62] ),
    .A1(_05544_),
    .S(_05417_),
    .X(_00283_));
 sky130_fd_sc_hd__mux2_1 _08463_ (.A0(mem_rdata[63]),
    .A1(cpu_wdata[63]),
    .S(cpu_write),
    .X(_05545_));
 sky130_fd_sc_hd__and2_2 _08464_ (.A(_05418_),
    .B(_05545_),
    .X(_05546_));
 sky130_fd_sc_hd__mux2_1 _08465_ (.A0(\data_array.data0[0][63] ),
    .A1(_05546_),
    .S(_05417_),
    .X(_00284_));
 sky130_fd_sc_hd__nor2_2 _08466_ (.A(_03507_),
    .B(_03511_),
    .Y(_05547_));
 sky130_fd_sc_hd__nand2_2 _08467_ (.A(_05360_),
    .B(_05547_),
    .Y(_05548_));
 sky130_fd_sc_hd__a21o_2 _08468_ (.A1(_05360_),
    .A2(_05547_),
    .B1(\tag_array.valid1[10] ),
    .X(_00285_));
 sky130_fd_sc_hd__and2_2 _08469_ (.A(_05360_),
    .B(_05416_),
    .X(_05549_));
 sky130_fd_sc_hd__or2_2 _08470_ (.A(\tag_array.valid1[0] ),
    .B(_05549_),
    .X(_00286_));
 sky130_fd_sc_hd__nand2_2 _08471_ (.A(_03506_),
    .B(_03515_),
    .Y(_05550_));
 sky130_fd_sc_hd__nand2b_2 _08472_ (.A_N(_05550_),
    .B(_05360_),
    .Y(_05551_));
 sky130_fd_sc_hd__a31o_2 _08473_ (.A1(_03506_),
    .A2(_03515_),
    .A3(_05360_),
    .B1(\tag_array.valid1[11] ),
    .X(_00287_));
 sky130_fd_sc_hd__nand2_2 _08474_ (.A(_03510_),
    .B(_03522_),
    .Y(_05552_));
 sky130_fd_sc_hd__or2_2 _08475_ (.A(_05353_),
    .B(_05552_),
    .X(_05553_));
 sky130_fd_sc_hd__nor2_2 _08476_ (.A(cpu_write),
    .B(_03146_),
    .Y(_05554_));
 sky130_fd_sc_hd__or4_2 _08477_ (.A(_05353_),
    .B(_05360_),
    .C(_05552_),
    .D(_05554_),
    .X(_05555_));
 sky130_fd_sc_hd__nand2b_2 _08478_ (.A_N(\tag_array.valid0[14] ),
    .B(_05555_),
    .Y(_00288_));
 sky130_fd_sc_hd__nor2_2 _08479_ (.A(_03507_),
    .B(_03514_),
    .Y(_05556_));
 sky130_fd_sc_hd__and2_2 _08480_ (.A(_05360_),
    .B(_05556_),
    .X(_05557_));
 sky130_fd_sc_hd__or2_2 _08481_ (.A(\tag_array.valid1[8] ),
    .B(_05557_),
    .X(_00289_));
 sky130_fd_sc_hd__nand2_2 _08482_ (.A(_03508_),
    .B(_03522_),
    .Y(_05558_));
 sky130_fd_sc_hd__or2_2 _08483_ (.A(_05353_),
    .B(_05558_),
    .X(_05559_));
 sky130_fd_sc_hd__or4_2 _08484_ (.A(_05353_),
    .B(_05360_),
    .C(_05554_),
    .D(_05558_),
    .X(_05560_));
 sky130_fd_sc_hd__nand2b_2 _08485_ (.A_N(\tag_array.valid0[13] ),
    .B(_05560_),
    .Y(_00290_));
 sky130_fd_sc_hd__a31o_2 _08486_ (.A1(_03515_),
    .A2(_03526_),
    .A3(_05360_),
    .B1(\tag_array.valid1[7] ),
    .X(_00291_));
 sky130_fd_sc_hd__nor2_2 _08487_ (.A(_03514_),
    .B(_03523_),
    .Y(_05561_));
 sky130_fd_sc_hd__or3_2 _08488_ (.A(_03514_),
    .B(_03523_),
    .C(_05353_),
    .X(_05562_));
 sky130_fd_sc_hd__or4b_2 _08489_ (.A(_05353_),
    .B(_05360_),
    .C(_05554_),
    .D_N(_05561_),
    .X(_05563_));
 sky130_fd_sc_hd__nand2b_2 _08490_ (.A_N(\tag_array.valid0[12] ),
    .B(_05563_),
    .Y(_00292_));
 sky130_fd_sc_hd__or2_2 _08491_ (.A(_05353_),
    .B(_05550_),
    .X(_05564_));
 sky130_fd_sc_hd__or4_2 _08492_ (.A(_05353_),
    .B(_05360_),
    .C(_05550_),
    .D(_05554_),
    .X(_05565_));
 sky130_fd_sc_hd__nand2b_2 _08493_ (.A_N(\tag_array.valid0[11] ),
    .B(_05565_),
    .Y(_00293_));
 sky130_fd_sc_hd__or3_2 _08494_ (.A(_03507_),
    .B(_03511_),
    .C(_05353_),
    .X(_05566_));
 sky130_fd_sc_hd__or4b_2 _08495_ (.A(_05353_),
    .B(_05360_),
    .C(_05554_),
    .D_N(_05547_),
    .X(_05567_));
 sky130_fd_sc_hd__nand2b_2 _08496_ (.A_N(\tag_array.valid0[10] ),
    .B(_05567_),
    .Y(_00294_));
 sky130_fd_sc_hd__or3_2 _08497_ (.A(_03514_),
    .B(_03519_),
    .C(_05353_),
    .X(_05568_));
 sky130_fd_sc_hd__or4b_2 _08498_ (.A(_05353_),
    .B(_05360_),
    .C(_05554_),
    .D_N(_05416_),
    .X(_05569_));
 sky130_fd_sc_hd__nand2b_2 _08499_ (.A_N(\tag_array.valid0[0] ),
    .B(_05569_),
    .Y(_00295_));
 sky130_fd_sc_hd__or3_2 _08500_ (.A(_03507_),
    .B(_03514_),
    .C(_05353_),
    .X(_05570_));
 sky130_fd_sc_hd__or4b_2 _08501_ (.A(_05353_),
    .B(_05360_),
    .C(_05554_),
    .D_N(_05556_),
    .X(_05571_));
 sky130_fd_sc_hd__nand2b_2 _08502_ (.A_N(\tag_array.valid0[8] ),
    .B(_05571_),
    .Y(_00296_));
 sky130_fd_sc_hd__or2_2 _08503_ (.A(_05353_),
    .B(_05361_),
    .X(_05572_));
 sky130_fd_sc_hd__or4_2 _08504_ (.A(_05353_),
    .B(_05360_),
    .C(_05361_),
    .D(_05554_),
    .X(_05573_));
 sky130_fd_sc_hd__nand2b_2 _08505_ (.A_N(\tag_array.valid0[7] ),
    .B(_05573_),
    .Y(_00297_));
 sky130_fd_sc_hd__nor2_2 _08506_ (.A(_03511_),
    .B(_03527_),
    .Y(_05574_));
 sky130_fd_sc_hd__or3_2 _08507_ (.A(_03511_),
    .B(_03527_),
    .C(_05353_),
    .X(_05575_));
 sky130_fd_sc_hd__or4b_2 _08508_ (.A(_05353_),
    .B(_05360_),
    .C(_05554_),
    .D_N(_05574_),
    .X(_05576_));
 sky130_fd_sc_hd__nand2b_2 _08509_ (.A_N(\tag_array.valid0[6] ),
    .B(_05576_),
    .Y(_00298_));
 sky130_fd_sc_hd__nor2_2 _08510_ (.A(_03509_),
    .B(_03527_),
    .Y(_05577_));
 sky130_fd_sc_hd__or3_2 _08511_ (.A(_03509_),
    .B(_03527_),
    .C(_05353_),
    .X(_05578_));
 sky130_fd_sc_hd__or4b_2 _08512_ (.A(_05353_),
    .B(_05360_),
    .C(_05554_),
    .D_N(_05577_),
    .X(_05579_));
 sky130_fd_sc_hd__nand2b_2 _08513_ (.A_N(\tag_array.valid0[5] ),
    .B(_05579_),
    .Y(_00299_));
 sky130_fd_sc_hd__nor2_2 _08514_ (.A(_03514_),
    .B(_03527_),
    .Y(_05580_));
 sky130_fd_sc_hd__or3_2 _08515_ (.A(_03514_),
    .B(_03527_),
    .C(_05353_),
    .X(_05581_));
 sky130_fd_sc_hd__or4b_2 _08516_ (.A(_05353_),
    .B(_05360_),
    .C(_05554_),
    .D_N(_05580_),
    .X(_05582_));
 sky130_fd_sc_hd__nand2b_2 _08517_ (.A_N(\tag_array.valid0[4] ),
    .B(_05582_),
    .Y(_00300_));
 sky130_fd_sc_hd__nor2_2 _08518_ (.A(_03516_),
    .B(_03519_),
    .Y(_05583_));
 sky130_fd_sc_hd__or3_2 _08519_ (.A(_03516_),
    .B(_03519_),
    .C(_05353_),
    .X(_05584_));
 sky130_fd_sc_hd__or4b_2 _08520_ (.A(_05353_),
    .B(_05360_),
    .C(_05554_),
    .D_N(_05583_),
    .X(_05585_));
 sky130_fd_sc_hd__nand2b_2 _08521_ (.A_N(\tag_array.valid0[3] ),
    .B(_05585_),
    .Y(_00301_));
 sky130_fd_sc_hd__or4b_2 _08522_ (.A(_05353_),
    .B(_05360_),
    .C(_05554_),
    .D_N(_05352_),
    .X(_05586_));
 sky130_fd_sc_hd__nand2b_2 _08523_ (.A_N(\tag_array.valid0[2] ),
    .B(_05586_),
    .Y(_00302_));
 sky130_fd_sc_hd__nor2_2 _08524_ (.A(_03509_),
    .B(_03519_),
    .Y(_05587_));
 sky130_fd_sc_hd__or3_2 _08525_ (.A(_03509_),
    .B(_03519_),
    .C(_05353_),
    .X(_05588_));
 sky130_fd_sc_hd__or4b_2 _08526_ (.A(_05353_),
    .B(_05360_),
    .C(_05554_),
    .D_N(_05587_),
    .X(_05589_));
 sky130_fd_sc_hd__nand2b_2 _08527_ (.A_N(\tag_array.valid0[1] ),
    .B(_05589_),
    .Y(_00303_));
 sky130_fd_sc_hd__nor2_2 _08528_ (.A(_03507_),
    .B(_03509_),
    .Y(_05590_));
 sky130_fd_sc_hd__nand2_2 _08529_ (.A(_05360_),
    .B(_05590_),
    .Y(_05591_));
 sky130_fd_sc_hd__a21o_2 _08530_ (.A1(_05360_),
    .A2(_05590_),
    .B1(\tag_array.valid1[9] ),
    .X(_00304_));
 sky130_fd_sc_hd__nand2b_2 _08531_ (.A_N(_05552_),
    .B(_05360_),
    .Y(_05592_));
 sky130_fd_sc_hd__a31o_2 _08532_ (.A1(_03510_),
    .A2(_03522_),
    .A3(_05360_),
    .B1(\tag_array.valid1[14] ),
    .X(_00305_));
 sky130_fd_sc_hd__nand2b_2 _08533_ (.A_N(_05558_),
    .B(_05360_),
    .Y(_05593_));
 sky130_fd_sc_hd__a31o_2 _08534_ (.A1(_03508_),
    .A2(_03522_),
    .A3(_05360_),
    .B1(\tag_array.valid1[13] ),
    .X(_00306_));
 sky130_fd_sc_hd__nand2_2 _08535_ (.A(_05360_),
    .B(_05561_),
    .Y(_05594_));
 sky130_fd_sc_hd__a21o_2 _08536_ (.A1(_05360_),
    .A2(_05561_),
    .B1(\tag_array.valid1[12] ),
    .X(_00307_));
 sky130_fd_sc_hd__nand2_2 _08537_ (.A(_03515_),
    .B(_03522_),
    .Y(_05595_));
 sky130_fd_sc_hd__or2_2 _08538_ (.A(_05353_),
    .B(_05595_),
    .X(_05596_));
 sky130_fd_sc_hd__or4_2 _08539_ (.A(_05353_),
    .B(_05360_),
    .C(_05554_),
    .D(_05595_),
    .X(_05597_));
 sky130_fd_sc_hd__nand2b_2 _08540_ (.A_N(\tag_array.valid0[15] ),
    .B(_05597_),
    .Y(_00308_));
 sky130_fd_sc_hd__mux2_1 _08541_ (.A0(_05365_),
    .A1(\tag_array.tag1[9][0] ),
    .S(_05591_),
    .X(_00309_));
 sky130_fd_sc_hd__mux2_1 _08542_ (.A0(_05367_),
    .A1(\tag_array.tag1[9][1] ),
    .S(_05591_),
    .X(_00310_));
 sky130_fd_sc_hd__mux2_1 _08543_ (.A0(_05369_),
    .A1(\tag_array.tag1[9][2] ),
    .S(_05591_),
    .X(_00311_));
 sky130_fd_sc_hd__mux2_1 _08544_ (.A0(_05371_),
    .A1(\tag_array.tag1[9][3] ),
    .S(_05591_),
    .X(_00312_));
 sky130_fd_sc_hd__mux2_1 _08545_ (.A0(_05373_),
    .A1(\tag_array.tag1[9][4] ),
    .S(_05591_),
    .X(_00313_));
 sky130_fd_sc_hd__mux2_1 _08546_ (.A0(_05375_),
    .A1(\tag_array.tag1[9][5] ),
    .S(_05591_),
    .X(_00314_));
 sky130_fd_sc_hd__mux2_1 _08547_ (.A0(_05377_),
    .A1(\tag_array.tag1[9][6] ),
    .S(_05591_),
    .X(_00315_));
 sky130_fd_sc_hd__mux2_1 _08548_ (.A0(_05379_),
    .A1(\tag_array.tag1[9][7] ),
    .S(_05591_),
    .X(_00316_));
 sky130_fd_sc_hd__mux2_1 _08549_ (.A0(_05381_),
    .A1(\tag_array.tag1[9][8] ),
    .S(_05591_),
    .X(_00317_));
 sky130_fd_sc_hd__mux2_1 _08550_ (.A0(_05383_),
    .A1(\tag_array.tag1[9][9] ),
    .S(_05591_),
    .X(_00318_));
 sky130_fd_sc_hd__mux2_1 _08551_ (.A0(_05385_),
    .A1(\tag_array.tag1[9][10] ),
    .S(_05591_),
    .X(_00319_));
 sky130_fd_sc_hd__mux2_1 _08552_ (.A0(_05387_),
    .A1(\tag_array.tag1[9][11] ),
    .S(_05591_),
    .X(_00320_));
 sky130_fd_sc_hd__mux2_1 _08553_ (.A0(_05389_),
    .A1(\tag_array.tag1[9][12] ),
    .S(_05591_),
    .X(_00321_));
 sky130_fd_sc_hd__mux2_1 _08554_ (.A0(_05391_),
    .A1(\tag_array.tag1[9][13] ),
    .S(_05591_),
    .X(_00322_));
 sky130_fd_sc_hd__mux2_1 _08555_ (.A0(_05393_),
    .A1(\tag_array.tag1[9][14] ),
    .S(_05591_),
    .X(_00323_));
 sky130_fd_sc_hd__mux2_1 _08556_ (.A0(_05395_),
    .A1(\tag_array.tag1[9][15] ),
    .S(_05591_),
    .X(_00324_));
 sky130_fd_sc_hd__mux2_1 _08557_ (.A0(_05397_),
    .A1(\tag_array.tag1[9][16] ),
    .S(_05591_),
    .X(_00325_));
 sky130_fd_sc_hd__mux2_1 _08558_ (.A0(_05399_),
    .A1(\tag_array.tag1[9][17] ),
    .S(_05591_),
    .X(_00326_));
 sky130_fd_sc_hd__mux2_1 _08559_ (.A0(_05401_),
    .A1(\tag_array.tag1[9][18] ),
    .S(_05591_),
    .X(_00327_));
 sky130_fd_sc_hd__mux2_1 _08560_ (.A0(_05403_),
    .A1(\tag_array.tag1[9][19] ),
    .S(_05591_),
    .X(_00328_));
 sky130_fd_sc_hd__mux2_1 _08561_ (.A0(_05405_),
    .A1(\tag_array.tag1[9][20] ),
    .S(_05591_),
    .X(_00329_));
 sky130_fd_sc_hd__mux2_1 _08562_ (.A0(_05407_),
    .A1(\tag_array.tag1[9][21] ),
    .S(_05591_),
    .X(_00330_));
 sky130_fd_sc_hd__mux2_1 _08563_ (.A0(_05409_),
    .A1(\tag_array.tag1[9][22] ),
    .S(_05591_),
    .X(_00331_));
 sky130_fd_sc_hd__mux2_1 _08564_ (.A0(_05411_),
    .A1(\tag_array.tag1[9][23] ),
    .S(_05591_),
    .X(_00332_));
 sky130_fd_sc_hd__mux2_1 _08565_ (.A0(_05413_),
    .A1(\tag_array.tag1[9][24] ),
    .S(_05591_),
    .X(_00333_));
 sky130_fd_sc_hd__nand2_2 _08566_ (.A(_05360_),
    .B(_05574_),
    .Y(_05598_));
 sky130_fd_sc_hd__a21o_2 _08567_ (.A1(_05360_),
    .A2(_05574_),
    .B1(\tag_array.valid1[6] ),
    .X(_00334_));
 sky130_fd_sc_hd__nand2_2 _08568_ (.A(_05360_),
    .B(_05577_),
    .Y(_05599_));
 sky130_fd_sc_hd__a21o_2 _08569_ (.A1(_05360_),
    .A2(_05577_),
    .B1(\tag_array.valid1[5] ),
    .X(_00335_));
 sky130_fd_sc_hd__and2_2 _08570_ (.A(_05360_),
    .B(_05580_),
    .X(_05600_));
 sky130_fd_sc_hd__or2_2 _08571_ (.A(\tag_array.valid1[4] ),
    .B(_05600_),
    .X(_00336_));
 sky130_fd_sc_hd__nand2_2 _08572_ (.A(_05360_),
    .B(_05583_),
    .Y(_05601_));
 sky130_fd_sc_hd__a21o_2 _08573_ (.A1(_05360_),
    .A2(_05583_),
    .B1(\tag_array.valid1[3] ),
    .X(_00337_));
 sky130_fd_sc_hd__and2_2 _08574_ (.A(_05352_),
    .B(_05360_),
    .X(_05602_));
 sky130_fd_sc_hd__or2_2 _08575_ (.A(\tag_array.valid1[2] ),
    .B(_05602_),
    .X(_00338_));
 sky130_fd_sc_hd__and2_2 _08576_ (.A(_05360_),
    .B(_05587_),
    .X(_05603_));
 sky130_fd_sc_hd__or2_2 _08577_ (.A(\tag_array.valid1[1] ),
    .B(_05603_),
    .X(_00339_));
 sky130_fd_sc_hd__nand2b_2 _08578_ (.A_N(_05595_),
    .B(_05360_),
    .Y(_05604_));
 sky130_fd_sc_hd__a31o_2 _08579_ (.A1(_03515_),
    .A2(_03522_),
    .A3(_05360_),
    .B1(\tag_array.valid1[15] ),
    .X(_00340_));
 sky130_fd_sc_hd__or3_2 _08580_ (.A(_03507_),
    .B(_03509_),
    .C(_05353_),
    .X(_05605_));
 sky130_fd_sc_hd__or4b_2 _08581_ (.A(_05353_),
    .B(_05360_),
    .C(_05554_),
    .D_N(_05590_),
    .X(_05606_));
 sky130_fd_sc_hd__nand2b_2 _08582_ (.A_N(\tag_array.valid0[9] ),
    .B(_05606_),
    .Y(_00341_));
 sky130_fd_sc_hd__mux2_1 _08583_ (.A0(_05365_),
    .A1(\tag_array.tag1[6][0] ),
    .S(_05598_),
    .X(_00342_));
 sky130_fd_sc_hd__mux2_1 _08584_ (.A0(_05367_),
    .A1(\tag_array.tag1[6][1] ),
    .S(_05598_),
    .X(_00343_));
 sky130_fd_sc_hd__mux2_1 _08585_ (.A0(_05369_),
    .A1(\tag_array.tag1[6][2] ),
    .S(_05598_),
    .X(_00344_));
 sky130_fd_sc_hd__mux2_1 _08586_ (.A0(_05371_),
    .A1(\tag_array.tag1[6][3] ),
    .S(_05598_),
    .X(_00345_));
 sky130_fd_sc_hd__mux2_1 _08587_ (.A0(_05373_),
    .A1(\tag_array.tag1[6][4] ),
    .S(_05598_),
    .X(_00346_));
 sky130_fd_sc_hd__mux2_1 _08588_ (.A0(_05375_),
    .A1(\tag_array.tag1[6][5] ),
    .S(_05598_),
    .X(_00347_));
 sky130_fd_sc_hd__mux2_1 _08589_ (.A0(_05377_),
    .A1(\tag_array.tag1[6][6] ),
    .S(_05598_),
    .X(_00348_));
 sky130_fd_sc_hd__mux2_1 _08590_ (.A0(_05379_),
    .A1(\tag_array.tag1[6][7] ),
    .S(_05598_),
    .X(_00349_));
 sky130_fd_sc_hd__mux2_1 _08591_ (.A0(_05381_),
    .A1(\tag_array.tag1[6][8] ),
    .S(_05598_),
    .X(_00350_));
 sky130_fd_sc_hd__mux2_1 _08592_ (.A0(_05383_),
    .A1(\tag_array.tag1[6][9] ),
    .S(_05598_),
    .X(_00351_));
 sky130_fd_sc_hd__mux2_1 _08593_ (.A0(_05385_),
    .A1(\tag_array.tag1[6][10] ),
    .S(_05598_),
    .X(_00352_));
 sky130_fd_sc_hd__mux2_1 _08594_ (.A0(_05387_),
    .A1(\tag_array.tag1[6][11] ),
    .S(_05598_),
    .X(_00353_));
 sky130_fd_sc_hd__mux2_1 _08595_ (.A0(_05389_),
    .A1(\tag_array.tag1[6][12] ),
    .S(_05598_),
    .X(_00354_));
 sky130_fd_sc_hd__mux2_1 _08596_ (.A0(_05391_),
    .A1(\tag_array.tag1[6][13] ),
    .S(_05598_),
    .X(_00355_));
 sky130_fd_sc_hd__mux2_1 _08597_ (.A0(_05393_),
    .A1(\tag_array.tag1[6][14] ),
    .S(_05598_),
    .X(_00356_));
 sky130_fd_sc_hd__mux2_1 _08598_ (.A0(_05395_),
    .A1(\tag_array.tag1[6][15] ),
    .S(_05598_),
    .X(_00357_));
 sky130_fd_sc_hd__mux2_1 _08599_ (.A0(_05397_),
    .A1(\tag_array.tag1[6][16] ),
    .S(_05598_),
    .X(_00358_));
 sky130_fd_sc_hd__mux2_1 _08600_ (.A0(_05399_),
    .A1(\tag_array.tag1[6][17] ),
    .S(_05598_),
    .X(_00359_));
 sky130_fd_sc_hd__mux2_1 _08601_ (.A0(_05401_),
    .A1(\tag_array.tag1[6][18] ),
    .S(_05598_),
    .X(_00360_));
 sky130_fd_sc_hd__mux2_1 _08602_ (.A0(_05403_),
    .A1(\tag_array.tag1[6][19] ),
    .S(_05598_),
    .X(_00361_));
 sky130_fd_sc_hd__mux2_1 _08603_ (.A0(_05405_),
    .A1(\tag_array.tag1[6][20] ),
    .S(_05598_),
    .X(_00362_));
 sky130_fd_sc_hd__mux2_1 _08604_ (.A0(_05407_),
    .A1(\tag_array.tag1[6][21] ),
    .S(_05598_),
    .X(_00363_));
 sky130_fd_sc_hd__mux2_1 _08605_ (.A0(_05409_),
    .A1(\tag_array.tag1[6][22] ),
    .S(_05598_),
    .X(_00364_));
 sky130_fd_sc_hd__mux2_1 _08606_ (.A0(_05411_),
    .A1(\tag_array.tag1[6][23] ),
    .S(_05598_),
    .X(_00365_));
 sky130_fd_sc_hd__mux2_1 _08607_ (.A0(_05413_),
    .A1(\tag_array.tag1[6][24] ),
    .S(_05598_),
    .X(_00366_));
 sky130_fd_sc_hd__mux2_1 _08608_ (.A0(_05365_),
    .A1(\tag_array.tag1[5][0] ),
    .S(_05599_),
    .X(_00367_));
 sky130_fd_sc_hd__mux2_1 _08609_ (.A0(_05367_),
    .A1(\tag_array.tag1[5][1] ),
    .S(_05599_),
    .X(_00368_));
 sky130_fd_sc_hd__mux2_1 _08610_ (.A0(_05369_),
    .A1(\tag_array.tag1[5][2] ),
    .S(_05599_),
    .X(_00369_));
 sky130_fd_sc_hd__mux2_1 _08611_ (.A0(_05371_),
    .A1(\tag_array.tag1[5][3] ),
    .S(_05599_),
    .X(_00370_));
 sky130_fd_sc_hd__mux2_1 _08612_ (.A0(_05373_),
    .A1(\tag_array.tag1[5][4] ),
    .S(_05599_),
    .X(_00371_));
 sky130_fd_sc_hd__mux2_1 _08613_ (.A0(_05375_),
    .A1(\tag_array.tag1[5][5] ),
    .S(_05599_),
    .X(_00372_));
 sky130_fd_sc_hd__mux2_1 _08614_ (.A0(_05377_),
    .A1(\tag_array.tag1[5][6] ),
    .S(_05599_),
    .X(_00373_));
 sky130_fd_sc_hd__mux2_1 _08615_ (.A0(_05379_),
    .A1(\tag_array.tag1[5][7] ),
    .S(_05599_),
    .X(_00374_));
 sky130_fd_sc_hd__mux2_1 _08616_ (.A0(_05381_),
    .A1(\tag_array.tag1[5][8] ),
    .S(_05599_),
    .X(_00375_));
 sky130_fd_sc_hd__mux2_1 _08617_ (.A0(_05383_),
    .A1(\tag_array.tag1[5][9] ),
    .S(_05599_),
    .X(_00376_));
 sky130_fd_sc_hd__mux2_1 _08618_ (.A0(_05385_),
    .A1(\tag_array.tag1[5][10] ),
    .S(_05599_),
    .X(_00377_));
 sky130_fd_sc_hd__mux2_1 _08619_ (.A0(_05387_),
    .A1(\tag_array.tag1[5][11] ),
    .S(_05599_),
    .X(_00378_));
 sky130_fd_sc_hd__mux2_1 _08620_ (.A0(_05389_),
    .A1(\tag_array.tag1[5][12] ),
    .S(_05599_),
    .X(_00379_));
 sky130_fd_sc_hd__mux2_1 _08621_ (.A0(_05391_),
    .A1(\tag_array.tag1[5][13] ),
    .S(_05599_),
    .X(_00380_));
 sky130_fd_sc_hd__mux2_1 _08622_ (.A0(_05393_),
    .A1(\tag_array.tag1[5][14] ),
    .S(_05599_),
    .X(_00381_));
 sky130_fd_sc_hd__mux2_1 _08623_ (.A0(_05395_),
    .A1(\tag_array.tag1[5][15] ),
    .S(_05599_),
    .X(_00382_));
 sky130_fd_sc_hd__mux2_1 _08624_ (.A0(_05397_),
    .A1(\tag_array.tag1[5][16] ),
    .S(_05599_),
    .X(_00383_));
 sky130_fd_sc_hd__mux2_1 _08625_ (.A0(_05399_),
    .A1(\tag_array.tag1[5][17] ),
    .S(_05599_),
    .X(_00384_));
 sky130_fd_sc_hd__mux2_1 _08626_ (.A0(_05401_),
    .A1(\tag_array.tag1[5][18] ),
    .S(_05599_),
    .X(_00385_));
 sky130_fd_sc_hd__mux2_1 _08627_ (.A0(_05403_),
    .A1(\tag_array.tag1[5][19] ),
    .S(_05599_),
    .X(_00386_));
 sky130_fd_sc_hd__mux2_1 _08628_ (.A0(_05405_),
    .A1(\tag_array.tag1[5][20] ),
    .S(_05599_),
    .X(_00387_));
 sky130_fd_sc_hd__mux2_1 _08629_ (.A0(_05407_),
    .A1(\tag_array.tag1[5][21] ),
    .S(_05599_),
    .X(_00388_));
 sky130_fd_sc_hd__mux2_1 _08630_ (.A0(_05409_),
    .A1(\tag_array.tag1[5][22] ),
    .S(_05599_),
    .X(_00389_));
 sky130_fd_sc_hd__mux2_1 _08631_ (.A0(_05411_),
    .A1(\tag_array.tag1[5][23] ),
    .S(_05599_),
    .X(_00390_));
 sky130_fd_sc_hd__mux2_1 _08632_ (.A0(_05413_),
    .A1(\tag_array.tag1[5][24] ),
    .S(_05599_),
    .X(_00391_));
 sky130_fd_sc_hd__mux2_1 _08633_ (.A0(\tag_array.tag1[4][0] ),
    .A1(_05365_),
    .S(_05600_),
    .X(_00392_));
 sky130_fd_sc_hd__mux2_1 _08634_ (.A0(\tag_array.tag1[4][1] ),
    .A1(_05367_),
    .S(_05600_),
    .X(_00393_));
 sky130_fd_sc_hd__mux2_1 _08635_ (.A0(\tag_array.tag1[4][2] ),
    .A1(_05369_),
    .S(_05600_),
    .X(_00394_));
 sky130_fd_sc_hd__mux2_1 _08636_ (.A0(\tag_array.tag1[4][3] ),
    .A1(_05371_),
    .S(_05600_),
    .X(_00395_));
 sky130_fd_sc_hd__mux2_1 _08637_ (.A0(\tag_array.tag1[4][4] ),
    .A1(_05373_),
    .S(_05600_),
    .X(_00396_));
 sky130_fd_sc_hd__mux2_1 _08638_ (.A0(\tag_array.tag1[4][5] ),
    .A1(_05375_),
    .S(_05600_),
    .X(_00397_));
 sky130_fd_sc_hd__mux2_1 _08639_ (.A0(\tag_array.tag1[4][6] ),
    .A1(_05377_),
    .S(_05600_),
    .X(_00398_));
 sky130_fd_sc_hd__mux2_1 _08640_ (.A0(\tag_array.tag1[4][7] ),
    .A1(_05379_),
    .S(_05600_),
    .X(_00399_));
 sky130_fd_sc_hd__mux2_1 _08641_ (.A0(\tag_array.tag1[4][8] ),
    .A1(_05381_),
    .S(_05600_),
    .X(_00400_));
 sky130_fd_sc_hd__mux2_1 _08642_ (.A0(\tag_array.tag1[4][9] ),
    .A1(_05383_),
    .S(_05600_),
    .X(_00401_));
 sky130_fd_sc_hd__mux2_1 _08643_ (.A0(\tag_array.tag1[4][10] ),
    .A1(_05385_),
    .S(_05600_),
    .X(_00402_));
 sky130_fd_sc_hd__mux2_1 _08644_ (.A0(\tag_array.tag1[4][11] ),
    .A1(_05387_),
    .S(_05600_),
    .X(_00403_));
 sky130_fd_sc_hd__mux2_1 _08645_ (.A0(\tag_array.tag1[4][12] ),
    .A1(_05389_),
    .S(_05600_),
    .X(_00404_));
 sky130_fd_sc_hd__mux2_1 _08646_ (.A0(\tag_array.tag1[4][13] ),
    .A1(_05391_),
    .S(_05600_),
    .X(_00405_));
 sky130_fd_sc_hd__mux2_1 _08647_ (.A0(\tag_array.tag1[4][14] ),
    .A1(_05393_),
    .S(_05600_),
    .X(_00406_));
 sky130_fd_sc_hd__mux2_1 _08648_ (.A0(\tag_array.tag1[4][15] ),
    .A1(_05395_),
    .S(_05600_),
    .X(_00407_));
 sky130_fd_sc_hd__mux2_1 _08649_ (.A0(\tag_array.tag1[4][16] ),
    .A1(_05397_),
    .S(_05600_),
    .X(_00408_));
 sky130_fd_sc_hd__mux2_1 _08650_ (.A0(\tag_array.tag1[4][17] ),
    .A1(_05399_),
    .S(_05600_),
    .X(_00409_));
 sky130_fd_sc_hd__mux2_1 _08651_ (.A0(\tag_array.tag1[4][18] ),
    .A1(_05401_),
    .S(_05600_),
    .X(_00410_));
 sky130_fd_sc_hd__mux2_1 _08652_ (.A0(\tag_array.tag1[4][19] ),
    .A1(_05403_),
    .S(_05600_),
    .X(_00411_));
 sky130_fd_sc_hd__mux2_1 _08653_ (.A0(\tag_array.tag1[4][20] ),
    .A1(_05405_),
    .S(_05600_),
    .X(_00412_));
 sky130_fd_sc_hd__mux2_1 _08654_ (.A0(\tag_array.tag1[4][21] ),
    .A1(_05407_),
    .S(_05600_),
    .X(_00413_));
 sky130_fd_sc_hd__mux2_1 _08655_ (.A0(\tag_array.tag1[4][22] ),
    .A1(_05409_),
    .S(_05600_),
    .X(_00414_));
 sky130_fd_sc_hd__mux2_1 _08656_ (.A0(\tag_array.tag1[4][23] ),
    .A1(_05411_),
    .S(_05600_),
    .X(_00415_));
 sky130_fd_sc_hd__mux2_1 _08657_ (.A0(\tag_array.tag1[4][24] ),
    .A1(_05413_),
    .S(_05600_),
    .X(_00416_));
 sky130_fd_sc_hd__mux2_1 _08658_ (.A0(_05365_),
    .A1(\tag_array.tag1[3][0] ),
    .S(_05601_),
    .X(_00417_));
 sky130_fd_sc_hd__mux2_1 _08659_ (.A0(_05367_),
    .A1(\tag_array.tag1[3][1] ),
    .S(_05601_),
    .X(_00418_));
 sky130_fd_sc_hd__mux2_1 _08660_ (.A0(_05369_),
    .A1(\tag_array.tag1[3][2] ),
    .S(_05601_),
    .X(_00419_));
 sky130_fd_sc_hd__mux2_1 _08661_ (.A0(_05371_),
    .A1(\tag_array.tag1[3][3] ),
    .S(_05601_),
    .X(_00420_));
 sky130_fd_sc_hd__mux2_1 _08662_ (.A0(_05373_),
    .A1(\tag_array.tag1[3][4] ),
    .S(_05601_),
    .X(_00421_));
 sky130_fd_sc_hd__mux2_1 _08663_ (.A0(_05375_),
    .A1(\tag_array.tag1[3][5] ),
    .S(_05601_),
    .X(_00422_));
 sky130_fd_sc_hd__mux2_1 _08664_ (.A0(_05377_),
    .A1(\tag_array.tag1[3][6] ),
    .S(_05601_),
    .X(_00423_));
 sky130_fd_sc_hd__mux2_1 _08665_ (.A0(_05379_),
    .A1(\tag_array.tag1[3][7] ),
    .S(_05601_),
    .X(_00424_));
 sky130_fd_sc_hd__mux2_1 _08666_ (.A0(_05381_),
    .A1(\tag_array.tag1[3][8] ),
    .S(_05601_),
    .X(_00425_));
 sky130_fd_sc_hd__mux2_1 _08667_ (.A0(_05383_),
    .A1(\tag_array.tag1[3][9] ),
    .S(_05601_),
    .X(_00426_));
 sky130_fd_sc_hd__mux2_1 _08668_ (.A0(_05385_),
    .A1(\tag_array.tag1[3][10] ),
    .S(_05601_),
    .X(_00427_));
 sky130_fd_sc_hd__mux2_1 _08669_ (.A0(_05387_),
    .A1(\tag_array.tag1[3][11] ),
    .S(_05601_),
    .X(_00428_));
 sky130_fd_sc_hd__mux2_1 _08670_ (.A0(_05389_),
    .A1(\tag_array.tag1[3][12] ),
    .S(_05601_),
    .X(_00429_));
 sky130_fd_sc_hd__mux2_1 _08671_ (.A0(_05391_),
    .A1(\tag_array.tag1[3][13] ),
    .S(_05601_),
    .X(_00430_));
 sky130_fd_sc_hd__mux2_1 _08672_ (.A0(_05393_),
    .A1(\tag_array.tag1[3][14] ),
    .S(_05601_),
    .X(_00431_));
 sky130_fd_sc_hd__mux2_1 _08673_ (.A0(_05395_),
    .A1(\tag_array.tag1[3][15] ),
    .S(_05601_),
    .X(_00432_));
 sky130_fd_sc_hd__mux2_1 _08674_ (.A0(_05397_),
    .A1(\tag_array.tag1[3][16] ),
    .S(_05601_),
    .X(_00433_));
 sky130_fd_sc_hd__mux2_1 _08675_ (.A0(_05399_),
    .A1(\tag_array.tag1[3][17] ),
    .S(_05601_),
    .X(_00434_));
 sky130_fd_sc_hd__mux2_1 _08676_ (.A0(_05401_),
    .A1(\tag_array.tag1[3][18] ),
    .S(_05601_),
    .X(_00435_));
 sky130_fd_sc_hd__mux2_1 _08677_ (.A0(_05403_),
    .A1(\tag_array.tag1[3][19] ),
    .S(_05601_),
    .X(_00436_));
 sky130_fd_sc_hd__mux2_1 _08678_ (.A0(_05405_),
    .A1(\tag_array.tag1[3][20] ),
    .S(_05601_),
    .X(_00437_));
 sky130_fd_sc_hd__mux2_1 _08679_ (.A0(_05407_),
    .A1(\tag_array.tag1[3][21] ),
    .S(_05601_),
    .X(_00438_));
 sky130_fd_sc_hd__mux2_1 _08680_ (.A0(_05409_),
    .A1(\tag_array.tag1[3][22] ),
    .S(_05601_),
    .X(_00439_));
 sky130_fd_sc_hd__mux2_1 _08681_ (.A0(_05411_),
    .A1(\tag_array.tag1[3][23] ),
    .S(_05601_),
    .X(_00440_));
 sky130_fd_sc_hd__mux2_1 _08682_ (.A0(_05413_),
    .A1(\tag_array.tag1[3][24] ),
    .S(_05601_),
    .X(_00441_));
 sky130_fd_sc_hd__mux2_1 _08683_ (.A0(\tag_array.tag1[2][0] ),
    .A1(_05365_),
    .S(_05602_),
    .X(_00442_));
 sky130_fd_sc_hd__mux2_1 _08684_ (.A0(\tag_array.tag1[2][1] ),
    .A1(_05367_),
    .S(_05602_),
    .X(_00443_));
 sky130_fd_sc_hd__mux2_1 _08685_ (.A0(\tag_array.tag1[2][2] ),
    .A1(_05369_),
    .S(_05602_),
    .X(_00444_));
 sky130_fd_sc_hd__mux2_1 _08686_ (.A0(\tag_array.tag1[2][3] ),
    .A1(_05371_),
    .S(_05602_),
    .X(_00445_));
 sky130_fd_sc_hd__mux2_1 _08687_ (.A0(\tag_array.tag1[2][4] ),
    .A1(_05373_),
    .S(_05602_),
    .X(_00446_));
 sky130_fd_sc_hd__mux2_1 _08688_ (.A0(\tag_array.tag1[2][5] ),
    .A1(_05375_),
    .S(_05602_),
    .X(_00447_));
 sky130_fd_sc_hd__mux2_1 _08689_ (.A0(\tag_array.tag1[2][6] ),
    .A1(_05377_),
    .S(_05602_),
    .X(_00448_));
 sky130_fd_sc_hd__mux2_1 _08690_ (.A0(\tag_array.tag1[2][7] ),
    .A1(_05379_),
    .S(_05602_),
    .X(_00449_));
 sky130_fd_sc_hd__mux2_1 _08691_ (.A0(\tag_array.tag1[2][8] ),
    .A1(_05381_),
    .S(_05602_),
    .X(_00450_));
 sky130_fd_sc_hd__mux2_1 _08692_ (.A0(\tag_array.tag1[2][9] ),
    .A1(_05383_),
    .S(_05602_),
    .X(_00451_));
 sky130_fd_sc_hd__mux2_1 _08693_ (.A0(\tag_array.tag1[2][10] ),
    .A1(_05385_),
    .S(_05602_),
    .X(_00452_));
 sky130_fd_sc_hd__mux2_1 _08694_ (.A0(\tag_array.tag1[2][11] ),
    .A1(_05387_),
    .S(_05602_),
    .X(_00453_));
 sky130_fd_sc_hd__mux2_1 _08695_ (.A0(\tag_array.tag1[2][12] ),
    .A1(_05389_),
    .S(_05602_),
    .X(_00454_));
 sky130_fd_sc_hd__mux2_1 _08696_ (.A0(\tag_array.tag1[2][13] ),
    .A1(_05391_),
    .S(_05602_),
    .X(_00455_));
 sky130_fd_sc_hd__mux2_1 _08697_ (.A0(\tag_array.tag1[2][14] ),
    .A1(_05393_),
    .S(_05602_),
    .X(_00456_));
 sky130_fd_sc_hd__mux2_1 _08698_ (.A0(\tag_array.tag1[2][15] ),
    .A1(_05395_),
    .S(_05602_),
    .X(_00457_));
 sky130_fd_sc_hd__mux2_1 _08699_ (.A0(\tag_array.tag1[2][16] ),
    .A1(_05397_),
    .S(_05602_),
    .X(_00458_));
 sky130_fd_sc_hd__mux2_1 _08700_ (.A0(\tag_array.tag1[2][17] ),
    .A1(_05399_),
    .S(_05602_),
    .X(_00459_));
 sky130_fd_sc_hd__mux2_1 _08701_ (.A0(\tag_array.tag1[2][18] ),
    .A1(_05401_),
    .S(_05602_),
    .X(_00460_));
 sky130_fd_sc_hd__mux2_1 _08702_ (.A0(\tag_array.tag1[2][19] ),
    .A1(_05403_),
    .S(_05602_),
    .X(_00461_));
 sky130_fd_sc_hd__mux2_1 _08703_ (.A0(\tag_array.tag1[2][20] ),
    .A1(_05405_),
    .S(_05602_),
    .X(_00462_));
 sky130_fd_sc_hd__mux2_1 _08704_ (.A0(\tag_array.tag1[2][21] ),
    .A1(_05407_),
    .S(_05602_),
    .X(_00463_));
 sky130_fd_sc_hd__mux2_1 _08705_ (.A0(\tag_array.tag1[2][22] ),
    .A1(_05409_),
    .S(_05602_),
    .X(_00464_));
 sky130_fd_sc_hd__mux2_1 _08706_ (.A0(\tag_array.tag1[2][23] ),
    .A1(_05411_),
    .S(_05602_),
    .X(_00465_));
 sky130_fd_sc_hd__mux2_1 _08707_ (.A0(\tag_array.tag1[2][24] ),
    .A1(_05413_),
    .S(_05602_),
    .X(_00466_));
 sky130_fd_sc_hd__mux2_1 _08708_ (.A0(\tag_array.tag1[1][0] ),
    .A1(_05365_),
    .S(_05603_),
    .X(_00467_));
 sky130_fd_sc_hd__mux2_1 _08709_ (.A0(\tag_array.tag1[1][1] ),
    .A1(_05367_),
    .S(_05603_),
    .X(_00468_));
 sky130_fd_sc_hd__mux2_1 _08710_ (.A0(\tag_array.tag1[1][2] ),
    .A1(_05369_),
    .S(_05603_),
    .X(_00469_));
 sky130_fd_sc_hd__mux2_1 _08711_ (.A0(\tag_array.tag1[1][3] ),
    .A1(_05371_),
    .S(_05603_),
    .X(_00470_));
 sky130_fd_sc_hd__mux2_1 _08712_ (.A0(\tag_array.tag1[1][4] ),
    .A1(_05373_),
    .S(_05603_),
    .X(_00471_));
 sky130_fd_sc_hd__mux2_1 _08713_ (.A0(\tag_array.tag1[1][5] ),
    .A1(_05375_),
    .S(_05603_),
    .X(_00472_));
 sky130_fd_sc_hd__mux2_1 _08714_ (.A0(\tag_array.tag1[1][6] ),
    .A1(_05377_),
    .S(_05603_),
    .X(_00473_));
 sky130_fd_sc_hd__mux2_1 _08715_ (.A0(\tag_array.tag1[1][7] ),
    .A1(_05379_),
    .S(_05603_),
    .X(_00474_));
 sky130_fd_sc_hd__mux2_1 _08716_ (.A0(\tag_array.tag1[1][8] ),
    .A1(_05381_),
    .S(_05603_),
    .X(_00475_));
 sky130_fd_sc_hd__mux2_1 _08717_ (.A0(\tag_array.tag1[1][9] ),
    .A1(_05383_),
    .S(_05603_),
    .X(_00476_));
 sky130_fd_sc_hd__mux2_1 _08718_ (.A0(\tag_array.tag1[1][10] ),
    .A1(_05385_),
    .S(_05603_),
    .X(_00477_));
 sky130_fd_sc_hd__mux2_1 _08719_ (.A0(\tag_array.tag1[1][11] ),
    .A1(_05387_),
    .S(_05603_),
    .X(_00478_));
 sky130_fd_sc_hd__mux2_1 _08720_ (.A0(\tag_array.tag1[1][12] ),
    .A1(_05389_),
    .S(_05603_),
    .X(_00479_));
 sky130_fd_sc_hd__mux2_1 _08721_ (.A0(\tag_array.tag1[1][13] ),
    .A1(_05391_),
    .S(_05603_),
    .X(_00480_));
 sky130_fd_sc_hd__mux2_1 _08722_ (.A0(\tag_array.tag1[1][14] ),
    .A1(_05393_),
    .S(_05603_),
    .X(_00481_));
 sky130_fd_sc_hd__mux2_1 _08723_ (.A0(\tag_array.tag1[1][15] ),
    .A1(_05395_),
    .S(_05603_),
    .X(_00482_));
 sky130_fd_sc_hd__mux2_1 _08724_ (.A0(\tag_array.tag1[1][16] ),
    .A1(_05397_),
    .S(_05603_),
    .X(_00483_));
 sky130_fd_sc_hd__mux2_1 _08725_ (.A0(\tag_array.tag1[1][17] ),
    .A1(_05399_),
    .S(_05603_),
    .X(_00484_));
 sky130_fd_sc_hd__mux2_1 _08726_ (.A0(\tag_array.tag1[1][18] ),
    .A1(_05401_),
    .S(_05603_),
    .X(_00485_));
 sky130_fd_sc_hd__mux2_1 _08727_ (.A0(\tag_array.tag1[1][19] ),
    .A1(_05403_),
    .S(_05603_),
    .X(_00486_));
 sky130_fd_sc_hd__mux2_1 _08728_ (.A0(\tag_array.tag1[1][20] ),
    .A1(_05405_),
    .S(_05603_),
    .X(_00487_));
 sky130_fd_sc_hd__mux2_1 _08729_ (.A0(\tag_array.tag1[1][21] ),
    .A1(_05407_),
    .S(_05603_),
    .X(_00488_));
 sky130_fd_sc_hd__mux2_1 _08730_ (.A0(\tag_array.tag1[1][22] ),
    .A1(_05409_),
    .S(_05603_),
    .X(_00489_));
 sky130_fd_sc_hd__mux2_1 _08731_ (.A0(\tag_array.tag1[1][23] ),
    .A1(_05411_),
    .S(_05603_),
    .X(_00490_));
 sky130_fd_sc_hd__mux2_1 _08732_ (.A0(\tag_array.tag1[1][24] ),
    .A1(_05413_),
    .S(_05603_),
    .X(_00491_));
 sky130_fd_sc_hd__mux2_1 _08733_ (.A0(_05365_),
    .A1(\tag_array.tag1[15][0] ),
    .S(_05604_),
    .X(_00492_));
 sky130_fd_sc_hd__mux2_1 _08734_ (.A0(_05367_),
    .A1(\tag_array.tag1[15][1] ),
    .S(_05604_),
    .X(_00493_));
 sky130_fd_sc_hd__mux2_1 _08735_ (.A0(_05369_),
    .A1(\tag_array.tag1[15][2] ),
    .S(_05604_),
    .X(_00494_));
 sky130_fd_sc_hd__mux2_1 _08736_ (.A0(_05371_),
    .A1(\tag_array.tag1[15][3] ),
    .S(_05604_),
    .X(_00495_));
 sky130_fd_sc_hd__mux2_1 _08737_ (.A0(_05373_),
    .A1(\tag_array.tag1[15][4] ),
    .S(_05604_),
    .X(_00496_));
 sky130_fd_sc_hd__mux2_1 _08738_ (.A0(_05375_),
    .A1(\tag_array.tag1[15][5] ),
    .S(_05604_),
    .X(_00497_));
 sky130_fd_sc_hd__mux2_1 _08739_ (.A0(_05377_),
    .A1(\tag_array.tag1[15][6] ),
    .S(_05604_),
    .X(_00498_));
 sky130_fd_sc_hd__mux2_1 _08740_ (.A0(_05379_),
    .A1(\tag_array.tag1[15][7] ),
    .S(_05604_),
    .X(_00499_));
 sky130_fd_sc_hd__mux2_1 _08741_ (.A0(_05381_),
    .A1(\tag_array.tag1[15][8] ),
    .S(_05604_),
    .X(_00500_));
 sky130_fd_sc_hd__mux2_1 _08742_ (.A0(_05383_),
    .A1(\tag_array.tag1[15][9] ),
    .S(_05604_),
    .X(_00501_));
 sky130_fd_sc_hd__mux2_1 _08743_ (.A0(_05385_),
    .A1(\tag_array.tag1[15][10] ),
    .S(_05604_),
    .X(_00502_));
 sky130_fd_sc_hd__mux2_1 _08744_ (.A0(_05387_),
    .A1(\tag_array.tag1[15][11] ),
    .S(_05604_),
    .X(_00503_));
 sky130_fd_sc_hd__mux2_1 _08745_ (.A0(_05389_),
    .A1(\tag_array.tag1[15][12] ),
    .S(_05604_),
    .X(_00504_));
 sky130_fd_sc_hd__mux2_1 _08746_ (.A0(_05391_),
    .A1(\tag_array.tag1[15][13] ),
    .S(_05604_),
    .X(_00505_));
 sky130_fd_sc_hd__mux2_1 _08747_ (.A0(_05393_),
    .A1(\tag_array.tag1[15][14] ),
    .S(_05604_),
    .X(_00506_));
 sky130_fd_sc_hd__mux2_1 _08748_ (.A0(_05395_),
    .A1(\tag_array.tag1[15][15] ),
    .S(_05604_),
    .X(_00507_));
 sky130_fd_sc_hd__mux2_1 _08749_ (.A0(_05397_),
    .A1(\tag_array.tag1[15][16] ),
    .S(_05604_),
    .X(_00508_));
 sky130_fd_sc_hd__mux2_1 _08750_ (.A0(_05399_),
    .A1(\tag_array.tag1[15][17] ),
    .S(_05604_),
    .X(_00509_));
 sky130_fd_sc_hd__mux2_1 _08751_ (.A0(_05401_),
    .A1(\tag_array.tag1[15][18] ),
    .S(_05604_),
    .X(_00510_));
 sky130_fd_sc_hd__mux2_1 _08752_ (.A0(_05403_),
    .A1(\tag_array.tag1[15][19] ),
    .S(_05604_),
    .X(_00511_));
 sky130_fd_sc_hd__mux2_1 _08753_ (.A0(_05405_),
    .A1(\tag_array.tag1[15][20] ),
    .S(_05604_),
    .X(_00512_));
 sky130_fd_sc_hd__mux2_1 _08754_ (.A0(_05407_),
    .A1(\tag_array.tag1[15][21] ),
    .S(_05604_),
    .X(_00513_));
 sky130_fd_sc_hd__mux2_1 _08755_ (.A0(_05409_),
    .A1(\tag_array.tag1[15][22] ),
    .S(_05604_),
    .X(_00514_));
 sky130_fd_sc_hd__mux2_1 _08756_ (.A0(_05411_),
    .A1(\tag_array.tag1[15][23] ),
    .S(_05604_),
    .X(_00515_));
 sky130_fd_sc_hd__mux2_1 _08757_ (.A0(_05413_),
    .A1(\tag_array.tag1[15][24] ),
    .S(_05604_),
    .X(_00516_));
 sky130_fd_sc_hd__mux2_1 _08758_ (.A0(_05365_),
    .A1(\tag_array.tag0[9][0] ),
    .S(_05606_),
    .X(_00517_));
 sky130_fd_sc_hd__mux2_1 _08759_ (.A0(_05367_),
    .A1(\tag_array.tag0[9][1] ),
    .S(_05606_),
    .X(_00518_));
 sky130_fd_sc_hd__mux2_1 _08760_ (.A0(_05369_),
    .A1(\tag_array.tag0[9][2] ),
    .S(_05606_),
    .X(_00519_));
 sky130_fd_sc_hd__mux2_1 _08761_ (.A0(_05371_),
    .A1(\tag_array.tag0[9][3] ),
    .S(_05606_),
    .X(_00520_));
 sky130_fd_sc_hd__mux2_1 _08762_ (.A0(_05373_),
    .A1(\tag_array.tag0[9][4] ),
    .S(_05606_),
    .X(_00521_));
 sky130_fd_sc_hd__mux2_1 _08763_ (.A0(_05375_),
    .A1(\tag_array.tag0[9][5] ),
    .S(_05606_),
    .X(_00522_));
 sky130_fd_sc_hd__mux2_1 _08764_ (.A0(_05377_),
    .A1(\tag_array.tag0[9][6] ),
    .S(_05606_),
    .X(_00523_));
 sky130_fd_sc_hd__mux2_1 _08765_ (.A0(_05379_),
    .A1(\tag_array.tag0[9][7] ),
    .S(_05606_),
    .X(_00524_));
 sky130_fd_sc_hd__mux2_1 _08766_ (.A0(_05381_),
    .A1(\tag_array.tag0[9][8] ),
    .S(_05606_),
    .X(_00525_));
 sky130_fd_sc_hd__mux2_1 _08767_ (.A0(_05383_),
    .A1(\tag_array.tag0[9][9] ),
    .S(_05606_),
    .X(_00526_));
 sky130_fd_sc_hd__mux2_1 _08768_ (.A0(_05385_),
    .A1(\tag_array.tag0[9][10] ),
    .S(_05606_),
    .X(_00527_));
 sky130_fd_sc_hd__mux2_1 _08769_ (.A0(_05387_),
    .A1(\tag_array.tag0[9][11] ),
    .S(_05606_),
    .X(_00528_));
 sky130_fd_sc_hd__mux2_1 _08770_ (.A0(_05389_),
    .A1(\tag_array.tag0[9][12] ),
    .S(_05606_),
    .X(_00529_));
 sky130_fd_sc_hd__mux2_1 _08771_ (.A0(_05391_),
    .A1(\tag_array.tag0[9][13] ),
    .S(_05606_),
    .X(_00530_));
 sky130_fd_sc_hd__mux2_1 _08772_ (.A0(_05393_),
    .A1(\tag_array.tag0[9][14] ),
    .S(_05606_),
    .X(_00531_));
 sky130_fd_sc_hd__mux2_1 _08773_ (.A0(_05395_),
    .A1(\tag_array.tag0[9][15] ),
    .S(_05606_),
    .X(_00532_));
 sky130_fd_sc_hd__mux2_1 _08774_ (.A0(_05397_),
    .A1(\tag_array.tag0[9][16] ),
    .S(_05606_),
    .X(_00533_));
 sky130_fd_sc_hd__mux2_1 _08775_ (.A0(_05399_),
    .A1(\tag_array.tag0[9][17] ),
    .S(_05606_),
    .X(_00534_));
 sky130_fd_sc_hd__mux2_1 _08776_ (.A0(_05401_),
    .A1(\tag_array.tag0[9][18] ),
    .S(_05606_),
    .X(_00535_));
 sky130_fd_sc_hd__mux2_1 _08777_ (.A0(_05403_),
    .A1(\tag_array.tag0[9][19] ),
    .S(_05606_),
    .X(_00536_));
 sky130_fd_sc_hd__mux2_1 _08778_ (.A0(_05405_),
    .A1(\tag_array.tag0[9][20] ),
    .S(_05606_),
    .X(_00537_));
 sky130_fd_sc_hd__mux2_1 _08779_ (.A0(_05407_),
    .A1(\tag_array.tag0[9][21] ),
    .S(_05606_),
    .X(_00538_));
 sky130_fd_sc_hd__mux2_1 _08780_ (.A0(_05409_),
    .A1(\tag_array.tag0[9][22] ),
    .S(_05606_),
    .X(_00539_));
 sky130_fd_sc_hd__mux2_1 _08781_ (.A0(_05411_),
    .A1(\tag_array.tag0[9][23] ),
    .S(_05606_),
    .X(_00540_));
 sky130_fd_sc_hd__mux2_1 _08782_ (.A0(_05413_),
    .A1(\tag_array.tag0[9][24] ),
    .S(_05606_),
    .X(_00541_));
 sky130_fd_sc_hd__and2_2 _08783_ (.A(_05415_),
    .B(_05556_),
    .X(_05607_));
 sky130_fd_sc_hd__mux2_1 _08784_ (.A0(\data_array.data0[8][0] ),
    .A1(_05420_),
    .S(_05607_),
    .X(_00542_));
 sky130_fd_sc_hd__mux2_1 _08785_ (.A0(\data_array.data0[8][1] ),
    .A1(_05422_),
    .S(_05607_),
    .X(_00543_));
 sky130_fd_sc_hd__mux2_1 _08786_ (.A0(\data_array.data0[8][2] ),
    .A1(_05424_),
    .S(_05607_),
    .X(_00544_));
 sky130_fd_sc_hd__mux2_1 _08787_ (.A0(\data_array.data0[8][3] ),
    .A1(_05426_),
    .S(_05607_),
    .X(_00545_));
 sky130_fd_sc_hd__mux2_1 _08788_ (.A0(\data_array.data0[8][4] ),
    .A1(_05428_),
    .S(_05607_),
    .X(_00546_));
 sky130_fd_sc_hd__mux2_1 _08789_ (.A0(\data_array.data0[8][5] ),
    .A1(_05430_),
    .S(_05607_),
    .X(_00547_));
 sky130_fd_sc_hd__mux2_1 _08790_ (.A0(\data_array.data0[8][6] ),
    .A1(_05432_),
    .S(_05607_),
    .X(_00548_));
 sky130_fd_sc_hd__mux2_1 _08791_ (.A0(\data_array.data0[8][7] ),
    .A1(_05434_),
    .S(_05607_),
    .X(_00549_));
 sky130_fd_sc_hd__mux2_1 _08792_ (.A0(\data_array.data0[8][8] ),
    .A1(_05436_),
    .S(_05607_),
    .X(_00550_));
 sky130_fd_sc_hd__mux2_1 _08793_ (.A0(\data_array.data0[8][9] ),
    .A1(_05438_),
    .S(_05607_),
    .X(_00551_));
 sky130_fd_sc_hd__mux2_1 _08794_ (.A0(\data_array.data0[8][10] ),
    .A1(_05440_),
    .S(_05607_),
    .X(_00552_));
 sky130_fd_sc_hd__mux2_1 _08795_ (.A0(\data_array.data0[8][11] ),
    .A1(_05442_),
    .S(_05607_),
    .X(_00553_));
 sky130_fd_sc_hd__mux2_1 _08796_ (.A0(\data_array.data0[8][12] ),
    .A1(_05444_),
    .S(_05607_),
    .X(_00554_));
 sky130_fd_sc_hd__mux2_1 _08797_ (.A0(\data_array.data0[8][13] ),
    .A1(_05446_),
    .S(_05607_),
    .X(_00555_));
 sky130_fd_sc_hd__mux2_1 _08798_ (.A0(\data_array.data0[8][14] ),
    .A1(_05448_),
    .S(_05607_),
    .X(_00556_));
 sky130_fd_sc_hd__mux2_1 _08799_ (.A0(\data_array.data0[8][15] ),
    .A1(_05450_),
    .S(_05607_),
    .X(_00557_));
 sky130_fd_sc_hd__mux2_1 _08800_ (.A0(\data_array.data0[8][16] ),
    .A1(_05452_),
    .S(_05607_),
    .X(_00558_));
 sky130_fd_sc_hd__mux2_1 _08801_ (.A0(\data_array.data0[8][17] ),
    .A1(_05454_),
    .S(_05607_),
    .X(_00559_));
 sky130_fd_sc_hd__mux2_1 _08802_ (.A0(\data_array.data0[8][18] ),
    .A1(_05456_),
    .S(_05607_),
    .X(_00560_));
 sky130_fd_sc_hd__mux2_1 _08803_ (.A0(\data_array.data0[8][19] ),
    .A1(_05458_),
    .S(_05607_),
    .X(_00561_));
 sky130_fd_sc_hd__mux2_1 _08804_ (.A0(\data_array.data0[8][20] ),
    .A1(_05460_),
    .S(_05607_),
    .X(_00562_));
 sky130_fd_sc_hd__mux2_1 _08805_ (.A0(\data_array.data0[8][21] ),
    .A1(_05462_),
    .S(_05607_),
    .X(_00563_));
 sky130_fd_sc_hd__mux2_1 _08806_ (.A0(\data_array.data0[8][22] ),
    .A1(_05464_),
    .S(_05607_),
    .X(_00564_));
 sky130_fd_sc_hd__mux2_1 _08807_ (.A0(\data_array.data0[8][23] ),
    .A1(_05466_),
    .S(_05607_),
    .X(_00565_));
 sky130_fd_sc_hd__mux2_1 _08808_ (.A0(\data_array.data0[8][24] ),
    .A1(_05468_),
    .S(_05607_),
    .X(_00566_));
 sky130_fd_sc_hd__mux2_1 _08809_ (.A0(\data_array.data0[8][25] ),
    .A1(_05470_),
    .S(_05607_),
    .X(_00567_));
 sky130_fd_sc_hd__mux2_1 _08810_ (.A0(\data_array.data0[8][26] ),
    .A1(_05472_),
    .S(_05607_),
    .X(_00568_));
 sky130_fd_sc_hd__mux2_1 _08811_ (.A0(\data_array.data0[8][27] ),
    .A1(_05474_),
    .S(_05607_),
    .X(_00569_));
 sky130_fd_sc_hd__mux2_1 _08812_ (.A0(\data_array.data0[8][28] ),
    .A1(_05476_),
    .S(_05607_),
    .X(_00570_));
 sky130_fd_sc_hd__mux2_1 _08813_ (.A0(\data_array.data0[8][29] ),
    .A1(_05478_),
    .S(_05607_),
    .X(_00571_));
 sky130_fd_sc_hd__mux2_1 _08814_ (.A0(\data_array.data0[8][30] ),
    .A1(_05480_),
    .S(_05607_),
    .X(_00572_));
 sky130_fd_sc_hd__mux2_1 _08815_ (.A0(\data_array.data0[8][31] ),
    .A1(_05482_),
    .S(_05607_),
    .X(_00573_));
 sky130_fd_sc_hd__mux2_1 _08816_ (.A0(\data_array.data0[8][32] ),
    .A1(_05484_),
    .S(_05607_),
    .X(_00574_));
 sky130_fd_sc_hd__mux2_1 _08817_ (.A0(\data_array.data0[8][33] ),
    .A1(_05486_),
    .S(_05607_),
    .X(_00575_));
 sky130_fd_sc_hd__mux2_1 _08818_ (.A0(\data_array.data0[8][34] ),
    .A1(_05488_),
    .S(_05607_),
    .X(_00576_));
 sky130_fd_sc_hd__mux2_1 _08819_ (.A0(\data_array.data0[8][35] ),
    .A1(_05490_),
    .S(_05607_),
    .X(_00577_));
 sky130_fd_sc_hd__mux2_1 _08820_ (.A0(\data_array.data0[8][36] ),
    .A1(_05492_),
    .S(_05607_),
    .X(_00578_));
 sky130_fd_sc_hd__mux2_1 _08821_ (.A0(\data_array.data0[8][37] ),
    .A1(_05494_),
    .S(_05607_),
    .X(_00579_));
 sky130_fd_sc_hd__mux2_1 _08822_ (.A0(\data_array.data0[8][38] ),
    .A1(_05496_),
    .S(_05607_),
    .X(_00580_));
 sky130_fd_sc_hd__mux2_1 _08823_ (.A0(\data_array.data0[8][39] ),
    .A1(_05498_),
    .S(_05607_),
    .X(_00581_));
 sky130_fd_sc_hd__mux2_1 _08824_ (.A0(\data_array.data0[8][40] ),
    .A1(_05500_),
    .S(_05607_),
    .X(_00582_));
 sky130_fd_sc_hd__mux2_1 _08825_ (.A0(\data_array.data0[8][41] ),
    .A1(_05502_),
    .S(_05607_),
    .X(_00583_));
 sky130_fd_sc_hd__mux2_1 _08826_ (.A0(\data_array.data0[8][42] ),
    .A1(_05504_),
    .S(_05607_),
    .X(_00584_));
 sky130_fd_sc_hd__mux2_1 _08827_ (.A0(\data_array.data0[8][43] ),
    .A1(_05506_),
    .S(_05607_),
    .X(_00585_));
 sky130_fd_sc_hd__mux2_1 _08828_ (.A0(\data_array.data0[8][44] ),
    .A1(_05508_),
    .S(_05607_),
    .X(_00586_));
 sky130_fd_sc_hd__mux2_1 _08829_ (.A0(\data_array.data0[8][45] ),
    .A1(_05510_),
    .S(_05607_),
    .X(_00587_));
 sky130_fd_sc_hd__mux2_1 _08830_ (.A0(\data_array.data0[8][46] ),
    .A1(_05512_),
    .S(_05607_),
    .X(_00588_));
 sky130_fd_sc_hd__mux2_1 _08831_ (.A0(\data_array.data0[8][47] ),
    .A1(_05514_),
    .S(_05607_),
    .X(_00589_));
 sky130_fd_sc_hd__mux2_1 _08832_ (.A0(\data_array.data0[8][48] ),
    .A1(_05516_),
    .S(_05607_),
    .X(_00590_));
 sky130_fd_sc_hd__mux2_1 _08833_ (.A0(\data_array.data0[8][49] ),
    .A1(_05518_),
    .S(_05607_),
    .X(_00591_));
 sky130_fd_sc_hd__mux2_1 _08834_ (.A0(\data_array.data0[8][50] ),
    .A1(_05520_),
    .S(_05607_),
    .X(_00592_));
 sky130_fd_sc_hd__mux2_1 _08835_ (.A0(\data_array.data0[8][51] ),
    .A1(_05522_),
    .S(_05607_),
    .X(_00593_));
 sky130_fd_sc_hd__mux2_1 _08836_ (.A0(\data_array.data0[8][52] ),
    .A1(_05524_),
    .S(_05607_),
    .X(_00594_));
 sky130_fd_sc_hd__mux2_1 _08837_ (.A0(\data_array.data0[8][53] ),
    .A1(_05526_),
    .S(_05607_),
    .X(_00595_));
 sky130_fd_sc_hd__mux2_1 _08838_ (.A0(\data_array.data0[8][54] ),
    .A1(_05528_),
    .S(_05607_),
    .X(_00596_));
 sky130_fd_sc_hd__mux2_1 _08839_ (.A0(\data_array.data0[8][55] ),
    .A1(_05530_),
    .S(_05607_),
    .X(_00597_));
 sky130_fd_sc_hd__mux2_1 _08840_ (.A0(\data_array.data0[8][56] ),
    .A1(_05532_),
    .S(_05607_),
    .X(_00598_));
 sky130_fd_sc_hd__mux2_1 _08841_ (.A0(\data_array.data0[8][57] ),
    .A1(_05534_),
    .S(_05607_),
    .X(_00599_));
 sky130_fd_sc_hd__mux2_1 _08842_ (.A0(\data_array.data0[8][58] ),
    .A1(_05536_),
    .S(_05607_),
    .X(_00600_));
 sky130_fd_sc_hd__mux2_1 _08843_ (.A0(\data_array.data0[8][59] ),
    .A1(_05538_),
    .S(_05607_),
    .X(_00601_));
 sky130_fd_sc_hd__mux2_1 _08844_ (.A0(\data_array.data0[8][60] ),
    .A1(_05540_),
    .S(_05607_),
    .X(_00602_));
 sky130_fd_sc_hd__mux2_1 _08845_ (.A0(\data_array.data0[8][61] ),
    .A1(_05542_),
    .S(_05607_),
    .X(_00603_));
 sky130_fd_sc_hd__mux2_1 _08846_ (.A0(\data_array.data0[8][62] ),
    .A1(_05544_),
    .S(_05607_),
    .X(_00604_));
 sky130_fd_sc_hd__mux2_1 _08847_ (.A0(\data_array.data0[8][63] ),
    .A1(_05546_),
    .S(_05607_),
    .X(_00605_));
 sky130_fd_sc_hd__or2_2 _08848_ (.A(_05361_),
    .B(_05414_),
    .X(_05608_));
 sky130_fd_sc_hd__mux2_1 _08849_ (.A0(_05420_),
    .A1(\data_array.data0[7][0] ),
    .S(_05608_),
    .X(_00606_));
 sky130_fd_sc_hd__mux2_1 _08850_ (.A0(_05422_),
    .A1(\data_array.data0[7][1] ),
    .S(_05608_),
    .X(_00607_));
 sky130_fd_sc_hd__mux2_1 _08851_ (.A0(_05424_),
    .A1(\data_array.data0[7][2] ),
    .S(_05608_),
    .X(_00608_));
 sky130_fd_sc_hd__mux2_1 _08852_ (.A0(_05426_),
    .A1(\data_array.data0[7][3] ),
    .S(_05608_),
    .X(_00609_));
 sky130_fd_sc_hd__mux2_1 _08853_ (.A0(_05428_),
    .A1(\data_array.data0[7][4] ),
    .S(_05608_),
    .X(_00610_));
 sky130_fd_sc_hd__mux2_1 _08854_ (.A0(_05430_),
    .A1(\data_array.data0[7][5] ),
    .S(_05608_),
    .X(_00611_));
 sky130_fd_sc_hd__mux2_1 _08855_ (.A0(_05432_),
    .A1(\data_array.data0[7][6] ),
    .S(_05608_),
    .X(_00612_));
 sky130_fd_sc_hd__mux2_1 _08856_ (.A0(_05434_),
    .A1(\data_array.data0[7][7] ),
    .S(_05608_),
    .X(_00613_));
 sky130_fd_sc_hd__mux2_1 _08857_ (.A0(_05436_),
    .A1(\data_array.data0[7][8] ),
    .S(_05608_),
    .X(_00614_));
 sky130_fd_sc_hd__mux2_1 _08858_ (.A0(_05438_),
    .A1(\data_array.data0[7][9] ),
    .S(_05608_),
    .X(_00615_));
 sky130_fd_sc_hd__mux2_1 _08859_ (.A0(_05440_),
    .A1(\data_array.data0[7][10] ),
    .S(_05608_),
    .X(_00616_));
 sky130_fd_sc_hd__mux2_1 _08860_ (.A0(_05442_),
    .A1(\data_array.data0[7][11] ),
    .S(_05608_),
    .X(_00617_));
 sky130_fd_sc_hd__mux2_1 _08861_ (.A0(_05444_),
    .A1(\data_array.data0[7][12] ),
    .S(_05608_),
    .X(_00618_));
 sky130_fd_sc_hd__mux2_1 _08862_ (.A0(_05446_),
    .A1(\data_array.data0[7][13] ),
    .S(_05608_),
    .X(_00619_));
 sky130_fd_sc_hd__mux2_1 _08863_ (.A0(_05448_),
    .A1(\data_array.data0[7][14] ),
    .S(_05608_),
    .X(_00620_));
 sky130_fd_sc_hd__mux2_1 _08864_ (.A0(_05450_),
    .A1(\data_array.data0[7][15] ),
    .S(_05608_),
    .X(_00621_));
 sky130_fd_sc_hd__mux2_1 _08865_ (.A0(_05452_),
    .A1(\data_array.data0[7][16] ),
    .S(_05608_),
    .X(_00622_));
 sky130_fd_sc_hd__mux2_1 _08866_ (.A0(_05454_),
    .A1(\data_array.data0[7][17] ),
    .S(_05608_),
    .X(_00623_));
 sky130_fd_sc_hd__mux2_1 _08867_ (.A0(_05456_),
    .A1(\data_array.data0[7][18] ),
    .S(_05608_),
    .X(_00624_));
 sky130_fd_sc_hd__mux2_1 _08868_ (.A0(_05458_),
    .A1(\data_array.data0[7][19] ),
    .S(_05608_),
    .X(_00625_));
 sky130_fd_sc_hd__mux2_1 _08869_ (.A0(_05460_),
    .A1(\data_array.data0[7][20] ),
    .S(_05608_),
    .X(_00626_));
 sky130_fd_sc_hd__mux2_1 _08870_ (.A0(_05462_),
    .A1(\data_array.data0[7][21] ),
    .S(_05608_),
    .X(_00627_));
 sky130_fd_sc_hd__mux2_1 _08871_ (.A0(_05464_),
    .A1(\data_array.data0[7][22] ),
    .S(_05608_),
    .X(_00628_));
 sky130_fd_sc_hd__mux2_1 _08872_ (.A0(_05466_),
    .A1(\data_array.data0[7][23] ),
    .S(_05608_),
    .X(_00629_));
 sky130_fd_sc_hd__mux2_1 _08873_ (.A0(_05468_),
    .A1(\data_array.data0[7][24] ),
    .S(_05608_),
    .X(_00630_));
 sky130_fd_sc_hd__mux2_1 _08874_ (.A0(_05470_),
    .A1(\data_array.data0[7][25] ),
    .S(_05608_),
    .X(_00631_));
 sky130_fd_sc_hd__mux2_1 _08875_ (.A0(_05472_),
    .A1(\data_array.data0[7][26] ),
    .S(_05608_),
    .X(_00632_));
 sky130_fd_sc_hd__mux2_1 _08876_ (.A0(_05474_),
    .A1(\data_array.data0[7][27] ),
    .S(_05608_),
    .X(_00633_));
 sky130_fd_sc_hd__mux2_1 _08877_ (.A0(_05476_),
    .A1(\data_array.data0[7][28] ),
    .S(_05608_),
    .X(_00634_));
 sky130_fd_sc_hd__mux2_1 _08878_ (.A0(_05478_),
    .A1(\data_array.data0[7][29] ),
    .S(_05608_),
    .X(_00635_));
 sky130_fd_sc_hd__mux2_1 _08879_ (.A0(_05480_),
    .A1(\data_array.data0[7][30] ),
    .S(_05608_),
    .X(_00636_));
 sky130_fd_sc_hd__mux2_1 _08880_ (.A0(_05482_),
    .A1(\data_array.data0[7][31] ),
    .S(_05608_),
    .X(_00637_));
 sky130_fd_sc_hd__mux2_1 _08881_ (.A0(_05484_),
    .A1(\data_array.data0[7][32] ),
    .S(_05608_),
    .X(_00638_));
 sky130_fd_sc_hd__mux2_1 _08882_ (.A0(_05486_),
    .A1(\data_array.data0[7][33] ),
    .S(_05608_),
    .X(_00639_));
 sky130_fd_sc_hd__mux2_1 _08883_ (.A0(_05488_),
    .A1(\data_array.data0[7][34] ),
    .S(_05608_),
    .X(_00640_));
 sky130_fd_sc_hd__mux2_1 _08884_ (.A0(_05490_),
    .A1(\data_array.data0[7][35] ),
    .S(_05608_),
    .X(_00641_));
 sky130_fd_sc_hd__mux2_1 _08885_ (.A0(_05492_),
    .A1(\data_array.data0[7][36] ),
    .S(_05608_),
    .X(_00642_));
 sky130_fd_sc_hd__mux2_1 _08886_ (.A0(_05494_),
    .A1(\data_array.data0[7][37] ),
    .S(_05608_),
    .X(_00643_));
 sky130_fd_sc_hd__mux2_1 _08887_ (.A0(_05496_),
    .A1(\data_array.data0[7][38] ),
    .S(_05608_),
    .X(_00644_));
 sky130_fd_sc_hd__mux2_1 _08888_ (.A0(_05498_),
    .A1(\data_array.data0[7][39] ),
    .S(_05608_),
    .X(_00645_));
 sky130_fd_sc_hd__mux2_1 _08889_ (.A0(_05500_),
    .A1(\data_array.data0[7][40] ),
    .S(_05608_),
    .X(_00646_));
 sky130_fd_sc_hd__mux2_1 _08890_ (.A0(_05502_),
    .A1(\data_array.data0[7][41] ),
    .S(_05608_),
    .X(_00647_));
 sky130_fd_sc_hd__mux2_1 _08891_ (.A0(_05504_),
    .A1(\data_array.data0[7][42] ),
    .S(_05608_),
    .X(_00648_));
 sky130_fd_sc_hd__mux2_1 _08892_ (.A0(_05506_),
    .A1(\data_array.data0[7][43] ),
    .S(_05608_),
    .X(_00649_));
 sky130_fd_sc_hd__mux2_1 _08893_ (.A0(_05508_),
    .A1(\data_array.data0[7][44] ),
    .S(_05608_),
    .X(_00650_));
 sky130_fd_sc_hd__mux2_1 _08894_ (.A0(_05510_),
    .A1(\data_array.data0[7][45] ),
    .S(_05608_),
    .X(_00651_));
 sky130_fd_sc_hd__mux2_1 _08895_ (.A0(_05512_),
    .A1(\data_array.data0[7][46] ),
    .S(_05608_),
    .X(_00652_));
 sky130_fd_sc_hd__mux2_1 _08896_ (.A0(_05514_),
    .A1(\data_array.data0[7][47] ),
    .S(_05608_),
    .X(_00653_));
 sky130_fd_sc_hd__mux2_1 _08897_ (.A0(_05516_),
    .A1(\data_array.data0[7][48] ),
    .S(_05608_),
    .X(_00654_));
 sky130_fd_sc_hd__mux2_1 _08898_ (.A0(_05518_),
    .A1(\data_array.data0[7][49] ),
    .S(_05608_),
    .X(_00655_));
 sky130_fd_sc_hd__mux2_1 _08899_ (.A0(_05520_),
    .A1(\data_array.data0[7][50] ),
    .S(_05608_),
    .X(_00656_));
 sky130_fd_sc_hd__mux2_1 _08900_ (.A0(_05522_),
    .A1(\data_array.data0[7][51] ),
    .S(_05608_),
    .X(_00657_));
 sky130_fd_sc_hd__mux2_1 _08901_ (.A0(_05524_),
    .A1(\data_array.data0[7][52] ),
    .S(_05608_),
    .X(_00658_));
 sky130_fd_sc_hd__mux2_1 _08902_ (.A0(_05526_),
    .A1(\data_array.data0[7][53] ),
    .S(_05608_),
    .X(_00659_));
 sky130_fd_sc_hd__mux2_1 _08903_ (.A0(_05528_),
    .A1(\data_array.data0[7][54] ),
    .S(_05608_),
    .X(_00660_));
 sky130_fd_sc_hd__mux2_1 _08904_ (.A0(_05530_),
    .A1(\data_array.data0[7][55] ),
    .S(_05608_),
    .X(_00661_));
 sky130_fd_sc_hd__mux2_1 _08905_ (.A0(_05532_),
    .A1(\data_array.data0[7][56] ),
    .S(_05608_),
    .X(_00662_));
 sky130_fd_sc_hd__mux2_1 _08906_ (.A0(_05534_),
    .A1(\data_array.data0[7][57] ),
    .S(_05608_),
    .X(_00663_));
 sky130_fd_sc_hd__mux2_1 _08907_ (.A0(_05536_),
    .A1(\data_array.data0[7][58] ),
    .S(_05608_),
    .X(_00664_));
 sky130_fd_sc_hd__mux2_1 _08908_ (.A0(_05538_),
    .A1(\data_array.data0[7][59] ),
    .S(_05608_),
    .X(_00665_));
 sky130_fd_sc_hd__mux2_1 _08909_ (.A0(_05540_),
    .A1(\data_array.data0[7][60] ),
    .S(_05608_),
    .X(_00666_));
 sky130_fd_sc_hd__mux2_1 _08910_ (.A0(_05542_),
    .A1(\data_array.data0[7][61] ),
    .S(_05608_),
    .X(_00667_));
 sky130_fd_sc_hd__mux2_1 _08911_ (.A0(_05544_),
    .A1(\data_array.data0[7][62] ),
    .S(_05608_),
    .X(_00668_));
 sky130_fd_sc_hd__mux2_1 _08912_ (.A0(_05546_),
    .A1(\data_array.data0[7][63] ),
    .S(_05608_),
    .X(_00669_));
 sky130_fd_sc_hd__nand2_2 _08913_ (.A(_05415_),
    .B(_05577_),
    .Y(_05609_));
 sky130_fd_sc_hd__mux2_1 _08914_ (.A0(_05420_),
    .A1(\data_array.data0[5][0] ),
    .S(_05609_),
    .X(_00670_));
 sky130_fd_sc_hd__mux2_1 _08915_ (.A0(_05422_),
    .A1(\data_array.data0[5][1] ),
    .S(_05609_),
    .X(_00671_));
 sky130_fd_sc_hd__mux2_1 _08916_ (.A0(_05424_),
    .A1(\data_array.data0[5][2] ),
    .S(_05609_),
    .X(_00672_));
 sky130_fd_sc_hd__mux2_1 _08917_ (.A0(_05426_),
    .A1(\data_array.data0[5][3] ),
    .S(_05609_),
    .X(_00673_));
 sky130_fd_sc_hd__mux2_1 _08918_ (.A0(_05428_),
    .A1(\data_array.data0[5][4] ),
    .S(_05609_),
    .X(_00674_));
 sky130_fd_sc_hd__mux2_1 _08919_ (.A0(_05430_),
    .A1(\data_array.data0[5][5] ),
    .S(_05609_),
    .X(_00675_));
 sky130_fd_sc_hd__mux2_1 _08920_ (.A0(_05432_),
    .A1(\data_array.data0[5][6] ),
    .S(_05609_),
    .X(_00676_));
 sky130_fd_sc_hd__mux2_1 _08921_ (.A0(_05434_),
    .A1(\data_array.data0[5][7] ),
    .S(_05609_),
    .X(_00677_));
 sky130_fd_sc_hd__mux2_1 _08922_ (.A0(_05436_),
    .A1(\data_array.data0[5][8] ),
    .S(_05609_),
    .X(_00678_));
 sky130_fd_sc_hd__mux2_1 _08923_ (.A0(_05438_),
    .A1(\data_array.data0[5][9] ),
    .S(_05609_),
    .X(_00679_));
 sky130_fd_sc_hd__mux2_1 _08924_ (.A0(_05440_),
    .A1(\data_array.data0[5][10] ),
    .S(_05609_),
    .X(_00680_));
 sky130_fd_sc_hd__mux2_1 _08925_ (.A0(_05442_),
    .A1(\data_array.data0[5][11] ),
    .S(_05609_),
    .X(_00681_));
 sky130_fd_sc_hd__mux2_1 _08926_ (.A0(_05444_),
    .A1(\data_array.data0[5][12] ),
    .S(_05609_),
    .X(_00682_));
 sky130_fd_sc_hd__mux2_1 _08927_ (.A0(_05446_),
    .A1(\data_array.data0[5][13] ),
    .S(_05609_),
    .X(_00683_));
 sky130_fd_sc_hd__mux2_1 _08928_ (.A0(_05448_),
    .A1(\data_array.data0[5][14] ),
    .S(_05609_),
    .X(_00684_));
 sky130_fd_sc_hd__mux2_1 _08929_ (.A0(_05450_),
    .A1(\data_array.data0[5][15] ),
    .S(_05609_),
    .X(_00685_));
 sky130_fd_sc_hd__mux2_1 _08930_ (.A0(_05452_),
    .A1(\data_array.data0[5][16] ),
    .S(_05609_),
    .X(_00686_));
 sky130_fd_sc_hd__mux2_1 _08931_ (.A0(_05454_),
    .A1(\data_array.data0[5][17] ),
    .S(_05609_),
    .X(_00687_));
 sky130_fd_sc_hd__mux2_1 _08932_ (.A0(_05456_),
    .A1(\data_array.data0[5][18] ),
    .S(_05609_),
    .X(_00688_));
 sky130_fd_sc_hd__mux2_1 _08933_ (.A0(_05458_),
    .A1(\data_array.data0[5][19] ),
    .S(_05609_),
    .X(_00689_));
 sky130_fd_sc_hd__mux2_1 _08934_ (.A0(_05460_),
    .A1(\data_array.data0[5][20] ),
    .S(_05609_),
    .X(_00690_));
 sky130_fd_sc_hd__mux2_1 _08935_ (.A0(_05462_),
    .A1(\data_array.data0[5][21] ),
    .S(_05609_),
    .X(_00691_));
 sky130_fd_sc_hd__mux2_1 _08936_ (.A0(_05464_),
    .A1(\data_array.data0[5][22] ),
    .S(_05609_),
    .X(_00692_));
 sky130_fd_sc_hd__mux2_1 _08937_ (.A0(_05466_),
    .A1(\data_array.data0[5][23] ),
    .S(_05609_),
    .X(_00693_));
 sky130_fd_sc_hd__mux2_1 _08938_ (.A0(_05468_),
    .A1(\data_array.data0[5][24] ),
    .S(_05609_),
    .X(_00694_));
 sky130_fd_sc_hd__mux2_1 _08939_ (.A0(_05470_),
    .A1(\data_array.data0[5][25] ),
    .S(_05609_),
    .X(_00695_));
 sky130_fd_sc_hd__mux2_1 _08940_ (.A0(_05472_),
    .A1(\data_array.data0[5][26] ),
    .S(_05609_),
    .X(_00696_));
 sky130_fd_sc_hd__mux2_1 _08941_ (.A0(_05474_),
    .A1(\data_array.data0[5][27] ),
    .S(_05609_),
    .X(_00697_));
 sky130_fd_sc_hd__mux2_1 _08942_ (.A0(_05476_),
    .A1(\data_array.data0[5][28] ),
    .S(_05609_),
    .X(_00698_));
 sky130_fd_sc_hd__mux2_1 _08943_ (.A0(_05478_),
    .A1(\data_array.data0[5][29] ),
    .S(_05609_),
    .X(_00699_));
 sky130_fd_sc_hd__mux2_1 _08944_ (.A0(_05480_),
    .A1(\data_array.data0[5][30] ),
    .S(_05609_),
    .X(_00700_));
 sky130_fd_sc_hd__mux2_1 _08945_ (.A0(_05482_),
    .A1(\data_array.data0[5][31] ),
    .S(_05609_),
    .X(_00701_));
 sky130_fd_sc_hd__mux2_1 _08946_ (.A0(_05484_),
    .A1(\data_array.data0[5][32] ),
    .S(_05609_),
    .X(_00702_));
 sky130_fd_sc_hd__mux2_1 _08947_ (.A0(_05486_),
    .A1(\data_array.data0[5][33] ),
    .S(_05609_),
    .X(_00703_));
 sky130_fd_sc_hd__mux2_1 _08948_ (.A0(_05488_),
    .A1(\data_array.data0[5][34] ),
    .S(_05609_),
    .X(_00704_));
 sky130_fd_sc_hd__mux2_1 _08949_ (.A0(_05490_),
    .A1(\data_array.data0[5][35] ),
    .S(_05609_),
    .X(_00705_));
 sky130_fd_sc_hd__mux2_1 _08950_ (.A0(_05492_),
    .A1(\data_array.data0[5][36] ),
    .S(_05609_),
    .X(_00706_));
 sky130_fd_sc_hd__mux2_1 _08951_ (.A0(_05494_),
    .A1(\data_array.data0[5][37] ),
    .S(_05609_),
    .X(_00707_));
 sky130_fd_sc_hd__mux2_1 _08952_ (.A0(_05496_),
    .A1(\data_array.data0[5][38] ),
    .S(_05609_),
    .X(_00708_));
 sky130_fd_sc_hd__mux2_1 _08953_ (.A0(_05498_),
    .A1(\data_array.data0[5][39] ),
    .S(_05609_),
    .X(_00709_));
 sky130_fd_sc_hd__mux2_1 _08954_ (.A0(_05500_),
    .A1(\data_array.data0[5][40] ),
    .S(_05609_),
    .X(_00710_));
 sky130_fd_sc_hd__mux2_1 _08955_ (.A0(_05502_),
    .A1(\data_array.data0[5][41] ),
    .S(_05609_),
    .X(_00711_));
 sky130_fd_sc_hd__mux2_1 _08956_ (.A0(_05504_),
    .A1(\data_array.data0[5][42] ),
    .S(_05609_),
    .X(_00712_));
 sky130_fd_sc_hd__mux2_1 _08957_ (.A0(_05506_),
    .A1(\data_array.data0[5][43] ),
    .S(_05609_),
    .X(_00713_));
 sky130_fd_sc_hd__mux2_1 _08958_ (.A0(_05508_),
    .A1(\data_array.data0[5][44] ),
    .S(_05609_),
    .X(_00714_));
 sky130_fd_sc_hd__mux2_1 _08959_ (.A0(_05510_),
    .A1(\data_array.data0[5][45] ),
    .S(_05609_),
    .X(_00715_));
 sky130_fd_sc_hd__mux2_1 _08960_ (.A0(_05512_),
    .A1(\data_array.data0[5][46] ),
    .S(_05609_),
    .X(_00716_));
 sky130_fd_sc_hd__mux2_1 _08961_ (.A0(_05514_),
    .A1(\data_array.data0[5][47] ),
    .S(_05609_),
    .X(_00717_));
 sky130_fd_sc_hd__mux2_1 _08962_ (.A0(_05516_),
    .A1(\data_array.data0[5][48] ),
    .S(_05609_),
    .X(_00718_));
 sky130_fd_sc_hd__mux2_1 _08963_ (.A0(_05518_),
    .A1(\data_array.data0[5][49] ),
    .S(_05609_),
    .X(_00719_));
 sky130_fd_sc_hd__mux2_1 _08964_ (.A0(_05520_),
    .A1(\data_array.data0[5][50] ),
    .S(_05609_),
    .X(_00720_));
 sky130_fd_sc_hd__mux2_1 _08965_ (.A0(_05522_),
    .A1(\data_array.data0[5][51] ),
    .S(_05609_),
    .X(_00721_));
 sky130_fd_sc_hd__mux2_1 _08966_ (.A0(_05524_),
    .A1(\data_array.data0[5][52] ),
    .S(_05609_),
    .X(_00722_));
 sky130_fd_sc_hd__mux2_1 _08967_ (.A0(_05526_),
    .A1(\data_array.data0[5][53] ),
    .S(_05609_),
    .X(_00723_));
 sky130_fd_sc_hd__mux2_1 _08968_ (.A0(_05528_),
    .A1(\data_array.data0[5][54] ),
    .S(_05609_),
    .X(_00724_));
 sky130_fd_sc_hd__mux2_1 _08969_ (.A0(_05530_),
    .A1(\data_array.data0[5][55] ),
    .S(_05609_),
    .X(_00725_));
 sky130_fd_sc_hd__mux2_1 _08970_ (.A0(_05532_),
    .A1(\data_array.data0[5][56] ),
    .S(_05609_),
    .X(_00726_));
 sky130_fd_sc_hd__mux2_1 _08971_ (.A0(_05534_),
    .A1(\data_array.data0[5][57] ),
    .S(_05609_),
    .X(_00727_));
 sky130_fd_sc_hd__mux2_1 _08972_ (.A0(_05536_),
    .A1(\data_array.data0[5][58] ),
    .S(_05609_),
    .X(_00728_));
 sky130_fd_sc_hd__mux2_1 _08973_ (.A0(_05538_),
    .A1(\data_array.data0[5][59] ),
    .S(_05609_),
    .X(_00729_));
 sky130_fd_sc_hd__mux2_1 _08974_ (.A0(_05540_),
    .A1(\data_array.data0[5][60] ),
    .S(_05609_),
    .X(_00730_));
 sky130_fd_sc_hd__mux2_1 _08975_ (.A0(_05542_),
    .A1(\data_array.data0[5][61] ),
    .S(_05609_),
    .X(_00731_));
 sky130_fd_sc_hd__mux2_1 _08976_ (.A0(_05544_),
    .A1(\data_array.data0[5][62] ),
    .S(_05609_),
    .X(_00732_));
 sky130_fd_sc_hd__mux2_1 _08977_ (.A0(_05546_),
    .A1(\data_array.data0[5][63] ),
    .S(_05609_),
    .X(_00733_));
 sky130_fd_sc_hd__and2_2 _08978_ (.A(_05415_),
    .B(_05580_),
    .X(_05610_));
 sky130_fd_sc_hd__mux2_1 _08979_ (.A0(\data_array.data0[4][0] ),
    .A1(_05420_),
    .S(_05610_),
    .X(_00734_));
 sky130_fd_sc_hd__mux2_1 _08980_ (.A0(\data_array.data0[4][1] ),
    .A1(_05422_),
    .S(_05610_),
    .X(_00735_));
 sky130_fd_sc_hd__mux2_1 _08981_ (.A0(\data_array.data0[4][2] ),
    .A1(_05424_),
    .S(_05610_),
    .X(_00736_));
 sky130_fd_sc_hd__mux2_1 _08982_ (.A0(\data_array.data0[4][3] ),
    .A1(_05426_),
    .S(_05610_),
    .X(_00737_));
 sky130_fd_sc_hd__mux2_1 _08983_ (.A0(\data_array.data0[4][4] ),
    .A1(_05428_),
    .S(_05610_),
    .X(_00738_));
 sky130_fd_sc_hd__mux2_1 _08984_ (.A0(\data_array.data0[4][5] ),
    .A1(_05430_),
    .S(_05610_),
    .X(_00739_));
 sky130_fd_sc_hd__mux2_1 _08985_ (.A0(\data_array.data0[4][6] ),
    .A1(_05432_),
    .S(_05610_),
    .X(_00740_));
 sky130_fd_sc_hd__mux2_1 _08986_ (.A0(\data_array.data0[4][7] ),
    .A1(_05434_),
    .S(_05610_),
    .X(_00741_));
 sky130_fd_sc_hd__mux2_1 _08987_ (.A0(\data_array.data0[4][8] ),
    .A1(_05436_),
    .S(_05610_),
    .X(_00742_));
 sky130_fd_sc_hd__mux2_1 _08988_ (.A0(\data_array.data0[4][9] ),
    .A1(_05438_),
    .S(_05610_),
    .X(_00743_));
 sky130_fd_sc_hd__mux2_1 _08989_ (.A0(\data_array.data0[4][10] ),
    .A1(_05440_),
    .S(_05610_),
    .X(_00744_));
 sky130_fd_sc_hd__mux2_1 _08990_ (.A0(\data_array.data0[4][11] ),
    .A1(_05442_),
    .S(_05610_),
    .X(_00745_));
 sky130_fd_sc_hd__mux2_1 _08991_ (.A0(\data_array.data0[4][12] ),
    .A1(_05444_),
    .S(_05610_),
    .X(_00746_));
 sky130_fd_sc_hd__mux2_1 _08992_ (.A0(\data_array.data0[4][13] ),
    .A1(_05446_),
    .S(_05610_),
    .X(_00747_));
 sky130_fd_sc_hd__mux2_1 _08993_ (.A0(\data_array.data0[4][14] ),
    .A1(_05448_),
    .S(_05610_),
    .X(_00748_));
 sky130_fd_sc_hd__mux2_1 _08994_ (.A0(\data_array.data0[4][15] ),
    .A1(_05450_),
    .S(_05610_),
    .X(_00749_));
 sky130_fd_sc_hd__mux2_1 _08995_ (.A0(\data_array.data0[4][16] ),
    .A1(_05452_),
    .S(_05610_),
    .X(_00750_));
 sky130_fd_sc_hd__mux2_1 _08996_ (.A0(\data_array.data0[4][17] ),
    .A1(_05454_),
    .S(_05610_),
    .X(_00751_));
 sky130_fd_sc_hd__mux2_1 _08997_ (.A0(\data_array.data0[4][18] ),
    .A1(_05456_),
    .S(_05610_),
    .X(_00752_));
 sky130_fd_sc_hd__mux2_1 _08998_ (.A0(\data_array.data0[4][19] ),
    .A1(_05458_),
    .S(_05610_),
    .X(_00753_));
 sky130_fd_sc_hd__mux2_1 _08999_ (.A0(\data_array.data0[4][20] ),
    .A1(_05460_),
    .S(_05610_),
    .X(_00754_));
 sky130_fd_sc_hd__mux2_1 _09000_ (.A0(\data_array.data0[4][21] ),
    .A1(_05462_),
    .S(_05610_),
    .X(_00755_));
 sky130_fd_sc_hd__mux2_1 _09001_ (.A0(\data_array.data0[4][22] ),
    .A1(_05464_),
    .S(_05610_),
    .X(_00756_));
 sky130_fd_sc_hd__mux2_1 _09002_ (.A0(\data_array.data0[4][23] ),
    .A1(_05466_),
    .S(_05610_),
    .X(_00757_));
 sky130_fd_sc_hd__mux2_1 _09003_ (.A0(\data_array.data0[4][24] ),
    .A1(_05468_),
    .S(_05610_),
    .X(_00758_));
 sky130_fd_sc_hd__mux2_1 _09004_ (.A0(\data_array.data0[4][25] ),
    .A1(_05470_),
    .S(_05610_),
    .X(_00759_));
 sky130_fd_sc_hd__mux2_1 _09005_ (.A0(\data_array.data0[4][26] ),
    .A1(_05472_),
    .S(_05610_),
    .X(_00760_));
 sky130_fd_sc_hd__mux2_1 _09006_ (.A0(\data_array.data0[4][27] ),
    .A1(_05474_),
    .S(_05610_),
    .X(_00761_));
 sky130_fd_sc_hd__mux2_1 _09007_ (.A0(\data_array.data0[4][28] ),
    .A1(_05476_),
    .S(_05610_),
    .X(_00762_));
 sky130_fd_sc_hd__mux2_1 _09008_ (.A0(\data_array.data0[4][29] ),
    .A1(_05478_),
    .S(_05610_),
    .X(_00763_));
 sky130_fd_sc_hd__mux2_1 _09009_ (.A0(\data_array.data0[4][30] ),
    .A1(_05480_),
    .S(_05610_),
    .X(_00764_));
 sky130_fd_sc_hd__mux2_1 _09010_ (.A0(\data_array.data0[4][31] ),
    .A1(_05482_),
    .S(_05610_),
    .X(_00765_));
 sky130_fd_sc_hd__mux2_1 _09011_ (.A0(\data_array.data0[4][32] ),
    .A1(_05484_),
    .S(_05610_),
    .X(_00766_));
 sky130_fd_sc_hd__mux2_1 _09012_ (.A0(\data_array.data0[4][33] ),
    .A1(_05486_),
    .S(_05610_),
    .X(_00767_));
 sky130_fd_sc_hd__mux2_1 _09013_ (.A0(\data_array.data0[4][34] ),
    .A1(_05488_),
    .S(_05610_),
    .X(_00768_));
 sky130_fd_sc_hd__mux2_1 _09014_ (.A0(\data_array.data0[4][35] ),
    .A1(_05490_),
    .S(_05610_),
    .X(_00769_));
 sky130_fd_sc_hd__mux2_1 _09015_ (.A0(\data_array.data0[4][36] ),
    .A1(_05492_),
    .S(_05610_),
    .X(_00770_));
 sky130_fd_sc_hd__mux2_1 _09016_ (.A0(\data_array.data0[4][37] ),
    .A1(_05494_),
    .S(_05610_),
    .X(_00771_));
 sky130_fd_sc_hd__mux2_1 _09017_ (.A0(\data_array.data0[4][38] ),
    .A1(_05496_),
    .S(_05610_),
    .X(_00772_));
 sky130_fd_sc_hd__mux2_1 _09018_ (.A0(\data_array.data0[4][39] ),
    .A1(_05498_),
    .S(_05610_),
    .X(_00773_));
 sky130_fd_sc_hd__mux2_1 _09019_ (.A0(\data_array.data0[4][40] ),
    .A1(_05500_),
    .S(_05610_),
    .X(_00774_));
 sky130_fd_sc_hd__mux2_1 _09020_ (.A0(\data_array.data0[4][41] ),
    .A1(_05502_),
    .S(_05610_),
    .X(_00775_));
 sky130_fd_sc_hd__mux2_1 _09021_ (.A0(\data_array.data0[4][42] ),
    .A1(_05504_),
    .S(_05610_),
    .X(_00776_));
 sky130_fd_sc_hd__mux2_1 _09022_ (.A0(\data_array.data0[4][43] ),
    .A1(_05506_),
    .S(_05610_),
    .X(_00777_));
 sky130_fd_sc_hd__mux2_1 _09023_ (.A0(\data_array.data0[4][44] ),
    .A1(_05508_),
    .S(_05610_),
    .X(_00778_));
 sky130_fd_sc_hd__mux2_1 _09024_ (.A0(\data_array.data0[4][45] ),
    .A1(_05510_),
    .S(_05610_),
    .X(_00779_));
 sky130_fd_sc_hd__mux2_1 _09025_ (.A0(\data_array.data0[4][46] ),
    .A1(_05512_),
    .S(_05610_),
    .X(_00780_));
 sky130_fd_sc_hd__mux2_1 _09026_ (.A0(\data_array.data0[4][47] ),
    .A1(_05514_),
    .S(_05610_),
    .X(_00781_));
 sky130_fd_sc_hd__mux2_1 _09027_ (.A0(\data_array.data0[4][48] ),
    .A1(_05516_),
    .S(_05610_),
    .X(_00782_));
 sky130_fd_sc_hd__mux2_1 _09028_ (.A0(\data_array.data0[4][49] ),
    .A1(_05518_),
    .S(_05610_),
    .X(_00783_));
 sky130_fd_sc_hd__mux2_1 _09029_ (.A0(\data_array.data0[4][50] ),
    .A1(_05520_),
    .S(_05610_),
    .X(_00784_));
 sky130_fd_sc_hd__mux2_1 _09030_ (.A0(\data_array.data0[4][51] ),
    .A1(_05522_),
    .S(_05610_),
    .X(_00785_));
 sky130_fd_sc_hd__mux2_1 _09031_ (.A0(\data_array.data0[4][52] ),
    .A1(_05524_),
    .S(_05610_),
    .X(_00786_));
 sky130_fd_sc_hd__mux2_1 _09032_ (.A0(\data_array.data0[4][53] ),
    .A1(_05526_),
    .S(_05610_),
    .X(_00787_));
 sky130_fd_sc_hd__mux2_1 _09033_ (.A0(\data_array.data0[4][54] ),
    .A1(_05528_),
    .S(_05610_),
    .X(_00788_));
 sky130_fd_sc_hd__mux2_1 _09034_ (.A0(\data_array.data0[4][55] ),
    .A1(_05530_),
    .S(_05610_),
    .X(_00789_));
 sky130_fd_sc_hd__mux2_1 _09035_ (.A0(\data_array.data0[4][56] ),
    .A1(_05532_),
    .S(_05610_),
    .X(_00790_));
 sky130_fd_sc_hd__mux2_1 _09036_ (.A0(\data_array.data0[4][57] ),
    .A1(_05534_),
    .S(_05610_),
    .X(_00791_));
 sky130_fd_sc_hd__mux2_1 _09037_ (.A0(\data_array.data0[4][58] ),
    .A1(_05536_),
    .S(_05610_),
    .X(_00792_));
 sky130_fd_sc_hd__mux2_1 _09038_ (.A0(\data_array.data0[4][59] ),
    .A1(_05538_),
    .S(_05610_),
    .X(_00793_));
 sky130_fd_sc_hd__mux2_1 _09039_ (.A0(\data_array.data0[4][60] ),
    .A1(_05540_),
    .S(_05610_),
    .X(_00794_));
 sky130_fd_sc_hd__mux2_1 _09040_ (.A0(\data_array.data0[4][61] ),
    .A1(_05542_),
    .S(_05610_),
    .X(_00795_));
 sky130_fd_sc_hd__mux2_1 _09041_ (.A0(\data_array.data0[4][62] ),
    .A1(_05544_),
    .S(_05610_),
    .X(_00796_));
 sky130_fd_sc_hd__mux2_1 _09042_ (.A0(\data_array.data0[4][63] ),
    .A1(_05546_),
    .S(_05610_),
    .X(_00797_));
 sky130_fd_sc_hd__nand2_2 _09043_ (.A(_05415_),
    .B(_05574_),
    .Y(_05611_));
 sky130_fd_sc_hd__mux2_1 _09044_ (.A0(_05420_),
    .A1(\data_array.data0[6][0] ),
    .S(_05611_),
    .X(_00798_));
 sky130_fd_sc_hd__mux2_1 _09045_ (.A0(_05422_),
    .A1(\data_array.data0[6][1] ),
    .S(_05611_),
    .X(_00799_));
 sky130_fd_sc_hd__mux2_1 _09046_ (.A0(_05424_),
    .A1(\data_array.data0[6][2] ),
    .S(_05611_),
    .X(_00800_));
 sky130_fd_sc_hd__mux2_1 _09047_ (.A0(_05426_),
    .A1(\data_array.data0[6][3] ),
    .S(_05611_),
    .X(_00801_));
 sky130_fd_sc_hd__mux2_1 _09048_ (.A0(_05428_),
    .A1(\data_array.data0[6][4] ),
    .S(_05611_),
    .X(_00802_));
 sky130_fd_sc_hd__mux2_1 _09049_ (.A0(_05430_),
    .A1(\data_array.data0[6][5] ),
    .S(_05611_),
    .X(_00803_));
 sky130_fd_sc_hd__mux2_1 _09050_ (.A0(_05432_),
    .A1(\data_array.data0[6][6] ),
    .S(_05611_),
    .X(_00804_));
 sky130_fd_sc_hd__mux2_1 _09051_ (.A0(_05434_),
    .A1(\data_array.data0[6][7] ),
    .S(_05611_),
    .X(_00805_));
 sky130_fd_sc_hd__mux2_1 _09052_ (.A0(_05436_),
    .A1(\data_array.data0[6][8] ),
    .S(_05611_),
    .X(_00806_));
 sky130_fd_sc_hd__mux2_1 _09053_ (.A0(_05438_),
    .A1(\data_array.data0[6][9] ),
    .S(_05611_),
    .X(_00807_));
 sky130_fd_sc_hd__mux2_1 _09054_ (.A0(_05440_),
    .A1(\data_array.data0[6][10] ),
    .S(_05611_),
    .X(_00808_));
 sky130_fd_sc_hd__mux2_1 _09055_ (.A0(_05442_),
    .A1(\data_array.data0[6][11] ),
    .S(_05611_),
    .X(_00809_));
 sky130_fd_sc_hd__mux2_1 _09056_ (.A0(_05444_),
    .A1(\data_array.data0[6][12] ),
    .S(_05611_),
    .X(_00810_));
 sky130_fd_sc_hd__mux2_1 _09057_ (.A0(_05446_),
    .A1(\data_array.data0[6][13] ),
    .S(_05611_),
    .X(_00811_));
 sky130_fd_sc_hd__mux2_1 _09058_ (.A0(_05448_),
    .A1(\data_array.data0[6][14] ),
    .S(_05611_),
    .X(_00812_));
 sky130_fd_sc_hd__mux2_1 _09059_ (.A0(_05450_),
    .A1(\data_array.data0[6][15] ),
    .S(_05611_),
    .X(_00813_));
 sky130_fd_sc_hd__mux2_1 _09060_ (.A0(_05452_),
    .A1(\data_array.data0[6][16] ),
    .S(_05611_),
    .X(_00814_));
 sky130_fd_sc_hd__mux2_1 _09061_ (.A0(_05454_),
    .A1(\data_array.data0[6][17] ),
    .S(_05611_),
    .X(_00815_));
 sky130_fd_sc_hd__mux2_1 _09062_ (.A0(_05456_),
    .A1(\data_array.data0[6][18] ),
    .S(_05611_),
    .X(_00816_));
 sky130_fd_sc_hd__mux2_1 _09063_ (.A0(_05458_),
    .A1(\data_array.data0[6][19] ),
    .S(_05611_),
    .X(_00817_));
 sky130_fd_sc_hd__mux2_1 _09064_ (.A0(_05460_),
    .A1(\data_array.data0[6][20] ),
    .S(_05611_),
    .X(_00818_));
 sky130_fd_sc_hd__mux2_1 _09065_ (.A0(_05462_),
    .A1(\data_array.data0[6][21] ),
    .S(_05611_),
    .X(_00819_));
 sky130_fd_sc_hd__mux2_1 _09066_ (.A0(_05464_),
    .A1(\data_array.data0[6][22] ),
    .S(_05611_),
    .X(_00820_));
 sky130_fd_sc_hd__mux2_1 _09067_ (.A0(_05466_),
    .A1(\data_array.data0[6][23] ),
    .S(_05611_),
    .X(_00821_));
 sky130_fd_sc_hd__mux2_1 _09068_ (.A0(_05468_),
    .A1(\data_array.data0[6][24] ),
    .S(_05611_),
    .X(_00822_));
 sky130_fd_sc_hd__mux2_1 _09069_ (.A0(_05470_),
    .A1(\data_array.data0[6][25] ),
    .S(_05611_),
    .X(_00823_));
 sky130_fd_sc_hd__mux2_1 _09070_ (.A0(_05472_),
    .A1(\data_array.data0[6][26] ),
    .S(_05611_),
    .X(_00824_));
 sky130_fd_sc_hd__mux2_1 _09071_ (.A0(_05474_),
    .A1(\data_array.data0[6][27] ),
    .S(_05611_),
    .X(_00825_));
 sky130_fd_sc_hd__mux2_1 _09072_ (.A0(_05476_),
    .A1(\data_array.data0[6][28] ),
    .S(_05611_),
    .X(_00826_));
 sky130_fd_sc_hd__mux2_1 _09073_ (.A0(_05478_),
    .A1(\data_array.data0[6][29] ),
    .S(_05611_),
    .X(_00827_));
 sky130_fd_sc_hd__mux2_1 _09074_ (.A0(_05480_),
    .A1(\data_array.data0[6][30] ),
    .S(_05611_),
    .X(_00828_));
 sky130_fd_sc_hd__mux2_1 _09075_ (.A0(_05482_),
    .A1(\data_array.data0[6][31] ),
    .S(_05611_),
    .X(_00829_));
 sky130_fd_sc_hd__mux2_1 _09076_ (.A0(_05484_),
    .A1(\data_array.data0[6][32] ),
    .S(_05611_),
    .X(_00830_));
 sky130_fd_sc_hd__mux2_1 _09077_ (.A0(_05486_),
    .A1(\data_array.data0[6][33] ),
    .S(_05611_),
    .X(_00831_));
 sky130_fd_sc_hd__mux2_1 _09078_ (.A0(_05488_),
    .A1(\data_array.data0[6][34] ),
    .S(_05611_),
    .X(_00832_));
 sky130_fd_sc_hd__mux2_1 _09079_ (.A0(_05490_),
    .A1(\data_array.data0[6][35] ),
    .S(_05611_),
    .X(_00833_));
 sky130_fd_sc_hd__mux2_1 _09080_ (.A0(_05492_),
    .A1(\data_array.data0[6][36] ),
    .S(_05611_),
    .X(_00834_));
 sky130_fd_sc_hd__mux2_1 _09081_ (.A0(_05494_),
    .A1(\data_array.data0[6][37] ),
    .S(_05611_),
    .X(_00835_));
 sky130_fd_sc_hd__mux2_1 _09082_ (.A0(_05496_),
    .A1(\data_array.data0[6][38] ),
    .S(_05611_),
    .X(_00836_));
 sky130_fd_sc_hd__mux2_1 _09083_ (.A0(_05498_),
    .A1(\data_array.data0[6][39] ),
    .S(_05611_),
    .X(_00837_));
 sky130_fd_sc_hd__mux2_1 _09084_ (.A0(_05500_),
    .A1(\data_array.data0[6][40] ),
    .S(_05611_),
    .X(_00838_));
 sky130_fd_sc_hd__mux2_1 _09085_ (.A0(_05502_),
    .A1(\data_array.data0[6][41] ),
    .S(_05611_),
    .X(_00839_));
 sky130_fd_sc_hd__mux2_1 _09086_ (.A0(_05504_),
    .A1(\data_array.data0[6][42] ),
    .S(_05611_),
    .X(_00840_));
 sky130_fd_sc_hd__mux2_1 _09087_ (.A0(_05506_),
    .A1(\data_array.data0[6][43] ),
    .S(_05611_),
    .X(_00841_));
 sky130_fd_sc_hd__mux2_1 _09088_ (.A0(_05508_),
    .A1(\data_array.data0[6][44] ),
    .S(_05611_),
    .X(_00842_));
 sky130_fd_sc_hd__mux2_1 _09089_ (.A0(_05510_),
    .A1(\data_array.data0[6][45] ),
    .S(_05611_),
    .X(_00843_));
 sky130_fd_sc_hd__mux2_1 _09090_ (.A0(_05512_),
    .A1(\data_array.data0[6][46] ),
    .S(_05611_),
    .X(_00844_));
 sky130_fd_sc_hd__mux2_1 _09091_ (.A0(_05514_),
    .A1(\data_array.data0[6][47] ),
    .S(_05611_),
    .X(_00845_));
 sky130_fd_sc_hd__mux2_1 _09092_ (.A0(_05516_),
    .A1(\data_array.data0[6][48] ),
    .S(_05611_),
    .X(_00846_));
 sky130_fd_sc_hd__mux2_1 _09093_ (.A0(_05518_),
    .A1(\data_array.data0[6][49] ),
    .S(_05611_),
    .X(_00847_));
 sky130_fd_sc_hd__mux2_1 _09094_ (.A0(_05520_),
    .A1(\data_array.data0[6][50] ),
    .S(_05611_),
    .X(_00848_));
 sky130_fd_sc_hd__mux2_1 _09095_ (.A0(_05522_),
    .A1(\data_array.data0[6][51] ),
    .S(_05611_),
    .X(_00849_));
 sky130_fd_sc_hd__mux2_1 _09096_ (.A0(_05524_),
    .A1(\data_array.data0[6][52] ),
    .S(_05611_),
    .X(_00850_));
 sky130_fd_sc_hd__mux2_1 _09097_ (.A0(_05526_),
    .A1(\data_array.data0[6][53] ),
    .S(_05611_),
    .X(_00851_));
 sky130_fd_sc_hd__mux2_1 _09098_ (.A0(_05528_),
    .A1(\data_array.data0[6][54] ),
    .S(_05611_),
    .X(_00852_));
 sky130_fd_sc_hd__mux2_1 _09099_ (.A0(_05530_),
    .A1(\data_array.data0[6][55] ),
    .S(_05611_),
    .X(_00853_));
 sky130_fd_sc_hd__mux2_1 _09100_ (.A0(_05532_),
    .A1(\data_array.data0[6][56] ),
    .S(_05611_),
    .X(_00854_));
 sky130_fd_sc_hd__mux2_1 _09101_ (.A0(_05534_),
    .A1(\data_array.data0[6][57] ),
    .S(_05611_),
    .X(_00855_));
 sky130_fd_sc_hd__mux2_1 _09102_ (.A0(_05536_),
    .A1(\data_array.data0[6][58] ),
    .S(_05611_),
    .X(_00856_));
 sky130_fd_sc_hd__mux2_1 _09103_ (.A0(_05538_),
    .A1(\data_array.data0[6][59] ),
    .S(_05611_),
    .X(_00857_));
 sky130_fd_sc_hd__mux2_1 _09104_ (.A0(_05540_),
    .A1(\data_array.data0[6][60] ),
    .S(_05611_),
    .X(_00858_));
 sky130_fd_sc_hd__mux2_1 _09105_ (.A0(_05542_),
    .A1(\data_array.data0[6][61] ),
    .S(_05611_),
    .X(_00859_));
 sky130_fd_sc_hd__mux2_1 _09106_ (.A0(_05544_),
    .A1(\data_array.data0[6][62] ),
    .S(_05611_),
    .X(_00860_));
 sky130_fd_sc_hd__mux2_1 _09107_ (.A0(_05546_),
    .A1(\data_array.data0[6][63] ),
    .S(_05611_),
    .X(_00861_));
 sky130_fd_sc_hd__mux2_1 _09108_ (.A0(_05420_),
    .A1(\data_array.data1[14][0] ),
    .S(_05592_),
    .X(_00862_));
 sky130_fd_sc_hd__mux2_1 _09109_ (.A0(_05422_),
    .A1(\data_array.data1[14][1] ),
    .S(_05592_),
    .X(_00863_));
 sky130_fd_sc_hd__mux2_1 _09110_ (.A0(_05424_),
    .A1(\data_array.data1[14][2] ),
    .S(_05592_),
    .X(_00864_));
 sky130_fd_sc_hd__mux2_1 _09111_ (.A0(_05426_),
    .A1(\data_array.data1[14][3] ),
    .S(_05592_),
    .X(_00865_));
 sky130_fd_sc_hd__mux2_1 _09112_ (.A0(_05428_),
    .A1(\data_array.data1[14][4] ),
    .S(_05592_),
    .X(_00866_));
 sky130_fd_sc_hd__mux2_1 _09113_ (.A0(_05430_),
    .A1(\data_array.data1[14][5] ),
    .S(_05592_),
    .X(_00867_));
 sky130_fd_sc_hd__mux2_1 _09114_ (.A0(_05432_),
    .A1(\data_array.data1[14][6] ),
    .S(_05592_),
    .X(_00868_));
 sky130_fd_sc_hd__mux2_1 _09115_ (.A0(_05434_),
    .A1(\data_array.data1[14][7] ),
    .S(_05592_),
    .X(_00869_));
 sky130_fd_sc_hd__mux2_1 _09116_ (.A0(_05436_),
    .A1(\data_array.data1[14][8] ),
    .S(_05592_),
    .X(_00870_));
 sky130_fd_sc_hd__mux2_1 _09117_ (.A0(_05438_),
    .A1(\data_array.data1[14][9] ),
    .S(_05592_),
    .X(_00871_));
 sky130_fd_sc_hd__mux2_1 _09118_ (.A0(_05440_),
    .A1(\data_array.data1[14][10] ),
    .S(_05592_),
    .X(_00872_));
 sky130_fd_sc_hd__mux2_1 _09119_ (.A0(_05442_),
    .A1(\data_array.data1[14][11] ),
    .S(_05592_),
    .X(_00873_));
 sky130_fd_sc_hd__mux2_1 _09120_ (.A0(_05444_),
    .A1(\data_array.data1[14][12] ),
    .S(_05592_),
    .X(_00874_));
 sky130_fd_sc_hd__mux2_1 _09121_ (.A0(_05446_),
    .A1(\data_array.data1[14][13] ),
    .S(_05592_),
    .X(_00875_));
 sky130_fd_sc_hd__mux2_1 _09122_ (.A0(_05448_),
    .A1(\data_array.data1[14][14] ),
    .S(_05592_),
    .X(_00876_));
 sky130_fd_sc_hd__mux2_1 _09123_ (.A0(_05450_),
    .A1(\data_array.data1[14][15] ),
    .S(_05592_),
    .X(_00877_));
 sky130_fd_sc_hd__mux2_1 _09124_ (.A0(_05452_),
    .A1(\data_array.data1[14][16] ),
    .S(_05592_),
    .X(_00878_));
 sky130_fd_sc_hd__mux2_1 _09125_ (.A0(_05454_),
    .A1(\data_array.data1[14][17] ),
    .S(_05592_),
    .X(_00879_));
 sky130_fd_sc_hd__mux2_1 _09126_ (.A0(_05456_),
    .A1(\data_array.data1[14][18] ),
    .S(_05592_),
    .X(_00880_));
 sky130_fd_sc_hd__mux2_1 _09127_ (.A0(_05458_),
    .A1(\data_array.data1[14][19] ),
    .S(_05592_),
    .X(_00881_));
 sky130_fd_sc_hd__mux2_1 _09128_ (.A0(_05460_),
    .A1(\data_array.data1[14][20] ),
    .S(_05592_),
    .X(_00882_));
 sky130_fd_sc_hd__mux2_1 _09129_ (.A0(_05462_),
    .A1(\data_array.data1[14][21] ),
    .S(_05592_),
    .X(_00883_));
 sky130_fd_sc_hd__mux2_1 _09130_ (.A0(_05464_),
    .A1(\data_array.data1[14][22] ),
    .S(_05592_),
    .X(_00884_));
 sky130_fd_sc_hd__mux2_1 _09131_ (.A0(_05466_),
    .A1(\data_array.data1[14][23] ),
    .S(_05592_),
    .X(_00885_));
 sky130_fd_sc_hd__mux2_1 _09132_ (.A0(_05468_),
    .A1(\data_array.data1[14][24] ),
    .S(_05592_),
    .X(_00886_));
 sky130_fd_sc_hd__mux2_1 _09133_ (.A0(_05470_),
    .A1(\data_array.data1[14][25] ),
    .S(_05592_),
    .X(_00887_));
 sky130_fd_sc_hd__mux2_1 _09134_ (.A0(_05472_),
    .A1(\data_array.data1[14][26] ),
    .S(_05592_),
    .X(_00888_));
 sky130_fd_sc_hd__mux2_1 _09135_ (.A0(_05474_),
    .A1(\data_array.data1[14][27] ),
    .S(_05592_),
    .X(_00889_));
 sky130_fd_sc_hd__mux2_1 _09136_ (.A0(_05476_),
    .A1(\data_array.data1[14][28] ),
    .S(_05592_),
    .X(_00890_));
 sky130_fd_sc_hd__mux2_1 _09137_ (.A0(_05478_),
    .A1(\data_array.data1[14][29] ),
    .S(_05592_),
    .X(_00891_));
 sky130_fd_sc_hd__mux2_1 _09138_ (.A0(_05480_),
    .A1(\data_array.data1[14][30] ),
    .S(_05592_),
    .X(_00892_));
 sky130_fd_sc_hd__mux2_1 _09139_ (.A0(_05482_),
    .A1(\data_array.data1[14][31] ),
    .S(_05592_),
    .X(_00893_));
 sky130_fd_sc_hd__mux2_1 _09140_ (.A0(_05484_),
    .A1(\data_array.data1[14][32] ),
    .S(_05592_),
    .X(_00894_));
 sky130_fd_sc_hd__mux2_1 _09141_ (.A0(_05486_),
    .A1(\data_array.data1[14][33] ),
    .S(_05592_),
    .X(_00895_));
 sky130_fd_sc_hd__mux2_1 _09142_ (.A0(_05488_),
    .A1(\data_array.data1[14][34] ),
    .S(_05592_),
    .X(_00896_));
 sky130_fd_sc_hd__mux2_1 _09143_ (.A0(_05490_),
    .A1(\data_array.data1[14][35] ),
    .S(_05592_),
    .X(_00897_));
 sky130_fd_sc_hd__mux2_1 _09144_ (.A0(_05492_),
    .A1(\data_array.data1[14][36] ),
    .S(_05592_),
    .X(_00898_));
 sky130_fd_sc_hd__mux2_1 _09145_ (.A0(_05494_),
    .A1(\data_array.data1[14][37] ),
    .S(_05592_),
    .X(_00899_));
 sky130_fd_sc_hd__mux2_1 _09146_ (.A0(_05496_),
    .A1(\data_array.data1[14][38] ),
    .S(_05592_),
    .X(_00900_));
 sky130_fd_sc_hd__mux2_1 _09147_ (.A0(_05498_),
    .A1(\data_array.data1[14][39] ),
    .S(_05592_),
    .X(_00901_));
 sky130_fd_sc_hd__mux2_1 _09148_ (.A0(_05500_),
    .A1(\data_array.data1[14][40] ),
    .S(_05592_),
    .X(_00902_));
 sky130_fd_sc_hd__mux2_1 _09149_ (.A0(_05502_),
    .A1(\data_array.data1[14][41] ),
    .S(_05592_),
    .X(_00903_));
 sky130_fd_sc_hd__mux2_1 _09150_ (.A0(_05504_),
    .A1(\data_array.data1[14][42] ),
    .S(_05592_),
    .X(_00904_));
 sky130_fd_sc_hd__mux2_1 _09151_ (.A0(_05506_),
    .A1(\data_array.data1[14][43] ),
    .S(_05592_),
    .X(_00905_));
 sky130_fd_sc_hd__mux2_1 _09152_ (.A0(_05508_),
    .A1(\data_array.data1[14][44] ),
    .S(_05592_),
    .X(_00906_));
 sky130_fd_sc_hd__mux2_1 _09153_ (.A0(_05510_),
    .A1(\data_array.data1[14][45] ),
    .S(_05592_),
    .X(_00907_));
 sky130_fd_sc_hd__mux2_1 _09154_ (.A0(_05512_),
    .A1(\data_array.data1[14][46] ),
    .S(_05592_),
    .X(_00908_));
 sky130_fd_sc_hd__mux2_1 _09155_ (.A0(_05514_),
    .A1(\data_array.data1[14][47] ),
    .S(_05592_),
    .X(_00909_));
 sky130_fd_sc_hd__mux2_1 _09156_ (.A0(_05516_),
    .A1(\data_array.data1[14][48] ),
    .S(_05592_),
    .X(_00910_));
 sky130_fd_sc_hd__mux2_1 _09157_ (.A0(_05518_),
    .A1(\data_array.data1[14][49] ),
    .S(_05592_),
    .X(_00911_));
 sky130_fd_sc_hd__mux2_1 _09158_ (.A0(_05520_),
    .A1(\data_array.data1[14][50] ),
    .S(_05592_),
    .X(_00912_));
 sky130_fd_sc_hd__mux2_1 _09159_ (.A0(_05522_),
    .A1(\data_array.data1[14][51] ),
    .S(_05592_),
    .X(_00913_));
 sky130_fd_sc_hd__mux2_1 _09160_ (.A0(_05524_),
    .A1(\data_array.data1[14][52] ),
    .S(_05592_),
    .X(_00914_));
 sky130_fd_sc_hd__mux2_1 _09161_ (.A0(_05526_),
    .A1(\data_array.data1[14][53] ),
    .S(_05592_),
    .X(_00915_));
 sky130_fd_sc_hd__mux2_1 _09162_ (.A0(_05528_),
    .A1(\data_array.data1[14][54] ),
    .S(_05592_),
    .X(_00916_));
 sky130_fd_sc_hd__mux2_1 _09163_ (.A0(_05530_),
    .A1(\data_array.data1[14][55] ),
    .S(_05592_),
    .X(_00917_));
 sky130_fd_sc_hd__mux2_1 _09164_ (.A0(_05532_),
    .A1(\data_array.data1[14][56] ),
    .S(_05592_),
    .X(_00918_));
 sky130_fd_sc_hd__mux2_1 _09165_ (.A0(_05534_),
    .A1(\data_array.data1[14][57] ),
    .S(_05592_),
    .X(_00919_));
 sky130_fd_sc_hd__mux2_1 _09166_ (.A0(_05536_),
    .A1(\data_array.data1[14][58] ),
    .S(_05592_),
    .X(_00920_));
 sky130_fd_sc_hd__mux2_1 _09167_ (.A0(_05538_),
    .A1(\data_array.data1[14][59] ),
    .S(_05592_),
    .X(_00921_));
 sky130_fd_sc_hd__mux2_1 _09168_ (.A0(_05540_),
    .A1(\data_array.data1[14][60] ),
    .S(_05592_),
    .X(_00922_));
 sky130_fd_sc_hd__mux2_1 _09169_ (.A0(_05542_),
    .A1(\data_array.data1[14][61] ),
    .S(_05592_),
    .X(_00923_));
 sky130_fd_sc_hd__mux2_1 _09170_ (.A0(_05544_),
    .A1(\data_array.data1[14][62] ),
    .S(_05592_),
    .X(_00924_));
 sky130_fd_sc_hd__mux2_1 _09171_ (.A0(_05546_),
    .A1(\data_array.data1[14][63] ),
    .S(_05592_),
    .X(_00925_));
 sky130_fd_sc_hd__mux2_1 _09172_ (.A0(_05365_),
    .A1(\tag_array.tag0[12][0] ),
    .S(_05563_),
    .X(_00926_));
 sky130_fd_sc_hd__mux2_1 _09173_ (.A0(_05367_),
    .A1(\tag_array.tag0[12][1] ),
    .S(_05563_),
    .X(_00927_));
 sky130_fd_sc_hd__mux2_1 _09174_ (.A0(_05369_),
    .A1(\tag_array.tag0[12][2] ),
    .S(_05563_),
    .X(_00928_));
 sky130_fd_sc_hd__mux2_1 _09175_ (.A0(_05371_),
    .A1(\tag_array.tag0[12][3] ),
    .S(_05563_),
    .X(_00929_));
 sky130_fd_sc_hd__mux2_1 _09176_ (.A0(_05373_),
    .A1(\tag_array.tag0[12][4] ),
    .S(_05563_),
    .X(_00930_));
 sky130_fd_sc_hd__mux2_1 _09177_ (.A0(_05375_),
    .A1(\tag_array.tag0[12][5] ),
    .S(_05563_),
    .X(_00931_));
 sky130_fd_sc_hd__mux2_1 _09178_ (.A0(_05377_),
    .A1(\tag_array.tag0[12][6] ),
    .S(_05563_),
    .X(_00932_));
 sky130_fd_sc_hd__mux2_1 _09179_ (.A0(_05379_),
    .A1(\tag_array.tag0[12][7] ),
    .S(_05563_),
    .X(_00933_));
 sky130_fd_sc_hd__mux2_1 _09180_ (.A0(_05381_),
    .A1(\tag_array.tag0[12][8] ),
    .S(_05563_),
    .X(_00934_));
 sky130_fd_sc_hd__mux2_1 _09181_ (.A0(_05383_),
    .A1(\tag_array.tag0[12][9] ),
    .S(_05563_),
    .X(_00935_));
 sky130_fd_sc_hd__mux2_1 _09182_ (.A0(_05385_),
    .A1(\tag_array.tag0[12][10] ),
    .S(_05563_),
    .X(_00936_));
 sky130_fd_sc_hd__mux2_1 _09183_ (.A0(_05387_),
    .A1(\tag_array.tag0[12][11] ),
    .S(_05563_),
    .X(_00937_));
 sky130_fd_sc_hd__mux2_1 _09184_ (.A0(_05389_),
    .A1(\tag_array.tag0[12][12] ),
    .S(_05563_),
    .X(_00938_));
 sky130_fd_sc_hd__mux2_1 _09185_ (.A0(_05391_),
    .A1(\tag_array.tag0[12][13] ),
    .S(_05563_),
    .X(_00939_));
 sky130_fd_sc_hd__mux2_1 _09186_ (.A0(_05393_),
    .A1(\tag_array.tag0[12][14] ),
    .S(_05563_),
    .X(_00940_));
 sky130_fd_sc_hd__mux2_1 _09187_ (.A0(_05395_),
    .A1(\tag_array.tag0[12][15] ),
    .S(_05563_),
    .X(_00941_));
 sky130_fd_sc_hd__mux2_1 _09188_ (.A0(_05397_),
    .A1(\tag_array.tag0[12][16] ),
    .S(_05563_),
    .X(_00942_));
 sky130_fd_sc_hd__mux2_1 _09189_ (.A0(_05399_),
    .A1(\tag_array.tag0[12][17] ),
    .S(_05563_),
    .X(_00943_));
 sky130_fd_sc_hd__mux2_1 _09190_ (.A0(_05401_),
    .A1(\tag_array.tag0[12][18] ),
    .S(_05563_),
    .X(_00944_));
 sky130_fd_sc_hd__mux2_1 _09191_ (.A0(_05403_),
    .A1(\tag_array.tag0[12][19] ),
    .S(_05563_),
    .X(_00945_));
 sky130_fd_sc_hd__mux2_1 _09192_ (.A0(_05405_),
    .A1(\tag_array.tag0[12][20] ),
    .S(_05563_),
    .X(_00946_));
 sky130_fd_sc_hd__mux2_1 _09193_ (.A0(_05407_),
    .A1(\tag_array.tag0[12][21] ),
    .S(_05563_),
    .X(_00947_));
 sky130_fd_sc_hd__mux2_1 _09194_ (.A0(_05409_),
    .A1(\tag_array.tag0[12][22] ),
    .S(_05563_),
    .X(_00948_));
 sky130_fd_sc_hd__mux2_1 _09195_ (.A0(_05411_),
    .A1(\tag_array.tag0[12][23] ),
    .S(_05563_),
    .X(_00949_));
 sky130_fd_sc_hd__mux2_1 _09196_ (.A0(_05413_),
    .A1(\tag_array.tag0[12][24] ),
    .S(_05563_),
    .X(_00950_));
 sky130_fd_sc_hd__mux2_1 _09197_ (.A0(_05365_),
    .A1(\tag_array.tag0[13][0] ),
    .S(_05560_),
    .X(_00951_));
 sky130_fd_sc_hd__mux2_1 _09198_ (.A0(_05367_),
    .A1(\tag_array.tag0[13][1] ),
    .S(_05560_),
    .X(_00952_));
 sky130_fd_sc_hd__mux2_1 _09199_ (.A0(_05369_),
    .A1(\tag_array.tag0[13][2] ),
    .S(_05560_),
    .X(_00953_));
 sky130_fd_sc_hd__mux2_1 _09200_ (.A0(_05371_),
    .A1(\tag_array.tag0[13][3] ),
    .S(_05560_),
    .X(_00954_));
 sky130_fd_sc_hd__mux2_1 _09201_ (.A0(_05373_),
    .A1(\tag_array.tag0[13][4] ),
    .S(_05560_),
    .X(_00955_));
 sky130_fd_sc_hd__mux2_1 _09202_ (.A0(_05375_),
    .A1(\tag_array.tag0[13][5] ),
    .S(_05560_),
    .X(_00956_));
 sky130_fd_sc_hd__mux2_1 _09203_ (.A0(_05377_),
    .A1(\tag_array.tag0[13][6] ),
    .S(_05560_),
    .X(_00957_));
 sky130_fd_sc_hd__mux2_1 _09204_ (.A0(_05379_),
    .A1(\tag_array.tag0[13][7] ),
    .S(_05560_),
    .X(_00958_));
 sky130_fd_sc_hd__mux2_1 _09205_ (.A0(_05381_),
    .A1(\tag_array.tag0[13][8] ),
    .S(_05560_),
    .X(_00959_));
 sky130_fd_sc_hd__mux2_1 _09206_ (.A0(_05383_),
    .A1(\tag_array.tag0[13][9] ),
    .S(_05560_),
    .X(_00960_));
 sky130_fd_sc_hd__mux2_1 _09207_ (.A0(_05385_),
    .A1(\tag_array.tag0[13][10] ),
    .S(_05560_),
    .X(_00961_));
 sky130_fd_sc_hd__mux2_1 _09208_ (.A0(_05387_),
    .A1(\tag_array.tag0[13][11] ),
    .S(_05560_),
    .X(_00962_));
 sky130_fd_sc_hd__mux2_1 _09209_ (.A0(_05389_),
    .A1(\tag_array.tag0[13][12] ),
    .S(_05560_),
    .X(_00963_));
 sky130_fd_sc_hd__mux2_1 _09210_ (.A0(_05391_),
    .A1(\tag_array.tag0[13][13] ),
    .S(_05560_),
    .X(_00964_));
 sky130_fd_sc_hd__mux2_1 _09211_ (.A0(_05393_),
    .A1(\tag_array.tag0[13][14] ),
    .S(_05560_),
    .X(_00965_));
 sky130_fd_sc_hd__mux2_1 _09212_ (.A0(_05395_),
    .A1(\tag_array.tag0[13][15] ),
    .S(_05560_),
    .X(_00966_));
 sky130_fd_sc_hd__mux2_1 _09213_ (.A0(_05397_),
    .A1(\tag_array.tag0[13][16] ),
    .S(_05560_),
    .X(_00967_));
 sky130_fd_sc_hd__mux2_1 _09214_ (.A0(_05399_),
    .A1(\tag_array.tag0[13][17] ),
    .S(_05560_),
    .X(_00968_));
 sky130_fd_sc_hd__mux2_1 _09215_ (.A0(_05401_),
    .A1(\tag_array.tag0[13][18] ),
    .S(_05560_),
    .X(_00969_));
 sky130_fd_sc_hd__mux2_1 _09216_ (.A0(_05403_),
    .A1(\tag_array.tag0[13][19] ),
    .S(_05560_),
    .X(_00970_));
 sky130_fd_sc_hd__mux2_1 _09217_ (.A0(_05405_),
    .A1(\tag_array.tag0[13][20] ),
    .S(_05560_),
    .X(_00971_));
 sky130_fd_sc_hd__mux2_1 _09218_ (.A0(_05407_),
    .A1(\tag_array.tag0[13][21] ),
    .S(_05560_),
    .X(_00972_));
 sky130_fd_sc_hd__mux2_1 _09219_ (.A0(_05409_),
    .A1(\tag_array.tag0[13][22] ),
    .S(_05560_),
    .X(_00973_));
 sky130_fd_sc_hd__mux2_1 _09220_ (.A0(_05411_),
    .A1(\tag_array.tag0[13][23] ),
    .S(_05560_),
    .X(_00974_));
 sky130_fd_sc_hd__mux2_1 _09221_ (.A0(_05413_),
    .A1(\tag_array.tag0[13][24] ),
    .S(_05560_),
    .X(_00975_));
 sky130_fd_sc_hd__mux2_1 _09222_ (.A0(_05365_),
    .A1(\tag_array.tag0[14][0] ),
    .S(_05555_),
    .X(_00976_));
 sky130_fd_sc_hd__mux2_1 _09223_ (.A0(_05367_),
    .A1(\tag_array.tag0[14][1] ),
    .S(_05555_),
    .X(_00977_));
 sky130_fd_sc_hd__mux2_1 _09224_ (.A0(_05369_),
    .A1(\tag_array.tag0[14][2] ),
    .S(_05555_),
    .X(_00978_));
 sky130_fd_sc_hd__mux2_1 _09225_ (.A0(_05371_),
    .A1(\tag_array.tag0[14][3] ),
    .S(_05555_),
    .X(_00979_));
 sky130_fd_sc_hd__mux2_1 _09226_ (.A0(_05373_),
    .A1(\tag_array.tag0[14][4] ),
    .S(_05555_),
    .X(_00980_));
 sky130_fd_sc_hd__mux2_1 _09227_ (.A0(_05375_),
    .A1(\tag_array.tag0[14][5] ),
    .S(_05555_),
    .X(_00981_));
 sky130_fd_sc_hd__mux2_1 _09228_ (.A0(_05377_),
    .A1(\tag_array.tag0[14][6] ),
    .S(_05555_),
    .X(_00982_));
 sky130_fd_sc_hd__mux2_1 _09229_ (.A0(_05379_),
    .A1(\tag_array.tag0[14][7] ),
    .S(_05555_),
    .X(_00983_));
 sky130_fd_sc_hd__mux2_1 _09230_ (.A0(_05381_),
    .A1(\tag_array.tag0[14][8] ),
    .S(_05555_),
    .X(_00984_));
 sky130_fd_sc_hd__mux2_1 _09231_ (.A0(_05383_),
    .A1(\tag_array.tag0[14][9] ),
    .S(_05555_),
    .X(_00985_));
 sky130_fd_sc_hd__mux2_1 _09232_ (.A0(_05385_),
    .A1(\tag_array.tag0[14][10] ),
    .S(_05555_),
    .X(_00986_));
 sky130_fd_sc_hd__mux2_1 _09233_ (.A0(_05387_),
    .A1(\tag_array.tag0[14][11] ),
    .S(_05555_),
    .X(_00987_));
 sky130_fd_sc_hd__mux2_1 _09234_ (.A0(_05389_),
    .A1(\tag_array.tag0[14][12] ),
    .S(_05555_),
    .X(_00988_));
 sky130_fd_sc_hd__mux2_1 _09235_ (.A0(_05391_),
    .A1(\tag_array.tag0[14][13] ),
    .S(_05555_),
    .X(_00989_));
 sky130_fd_sc_hd__mux2_1 _09236_ (.A0(_05393_),
    .A1(\tag_array.tag0[14][14] ),
    .S(_05555_),
    .X(_00990_));
 sky130_fd_sc_hd__mux2_1 _09237_ (.A0(_05395_),
    .A1(\tag_array.tag0[14][15] ),
    .S(_05555_),
    .X(_00991_));
 sky130_fd_sc_hd__mux2_1 _09238_ (.A0(_05397_),
    .A1(\tag_array.tag0[14][16] ),
    .S(_05555_),
    .X(_00992_));
 sky130_fd_sc_hd__mux2_1 _09239_ (.A0(_05399_),
    .A1(\tag_array.tag0[14][17] ),
    .S(_05555_),
    .X(_00993_));
 sky130_fd_sc_hd__mux2_1 _09240_ (.A0(_05401_),
    .A1(\tag_array.tag0[14][18] ),
    .S(_05555_),
    .X(_00994_));
 sky130_fd_sc_hd__mux2_1 _09241_ (.A0(_05403_),
    .A1(\tag_array.tag0[14][19] ),
    .S(_05555_),
    .X(_00995_));
 sky130_fd_sc_hd__mux2_1 _09242_ (.A0(_05405_),
    .A1(\tag_array.tag0[14][20] ),
    .S(_05555_),
    .X(_00996_));
 sky130_fd_sc_hd__mux2_1 _09243_ (.A0(_05407_),
    .A1(\tag_array.tag0[14][21] ),
    .S(_05555_),
    .X(_00997_));
 sky130_fd_sc_hd__mux2_1 _09244_ (.A0(_05409_),
    .A1(\tag_array.tag0[14][22] ),
    .S(_05555_),
    .X(_00998_));
 sky130_fd_sc_hd__mux2_1 _09245_ (.A0(_05411_),
    .A1(\tag_array.tag0[14][23] ),
    .S(_05555_),
    .X(_00999_));
 sky130_fd_sc_hd__mux2_1 _09246_ (.A0(_05413_),
    .A1(\tag_array.tag0[14][24] ),
    .S(_05555_),
    .X(_01000_));
 sky130_fd_sc_hd__mux2_1 _09247_ (.A0(_05365_),
    .A1(\tag_array.tag1[14][0] ),
    .S(_05592_),
    .X(_01001_));
 sky130_fd_sc_hd__mux2_1 _09248_ (.A0(_05367_),
    .A1(\tag_array.tag1[14][1] ),
    .S(_05592_),
    .X(_01002_));
 sky130_fd_sc_hd__mux2_1 _09249_ (.A0(_05369_),
    .A1(\tag_array.tag1[14][2] ),
    .S(_05592_),
    .X(_01003_));
 sky130_fd_sc_hd__mux2_1 _09250_ (.A0(_05371_),
    .A1(\tag_array.tag1[14][3] ),
    .S(_05592_),
    .X(_01004_));
 sky130_fd_sc_hd__mux2_1 _09251_ (.A0(_05373_),
    .A1(\tag_array.tag1[14][4] ),
    .S(_05592_),
    .X(_01005_));
 sky130_fd_sc_hd__mux2_1 _09252_ (.A0(_05375_),
    .A1(\tag_array.tag1[14][5] ),
    .S(_05592_),
    .X(_01006_));
 sky130_fd_sc_hd__mux2_1 _09253_ (.A0(_05377_),
    .A1(\tag_array.tag1[14][6] ),
    .S(_05592_),
    .X(_01007_));
 sky130_fd_sc_hd__mux2_1 _09254_ (.A0(_05379_),
    .A1(\tag_array.tag1[14][7] ),
    .S(_05592_),
    .X(_01008_));
 sky130_fd_sc_hd__mux2_1 _09255_ (.A0(_05381_),
    .A1(\tag_array.tag1[14][8] ),
    .S(_05592_),
    .X(_01009_));
 sky130_fd_sc_hd__mux2_1 _09256_ (.A0(_05383_),
    .A1(\tag_array.tag1[14][9] ),
    .S(_05592_),
    .X(_01010_));
 sky130_fd_sc_hd__mux2_1 _09257_ (.A0(_05385_),
    .A1(\tag_array.tag1[14][10] ),
    .S(_05592_),
    .X(_01011_));
 sky130_fd_sc_hd__mux2_1 _09258_ (.A0(_05387_),
    .A1(\tag_array.tag1[14][11] ),
    .S(_05592_),
    .X(_01012_));
 sky130_fd_sc_hd__mux2_1 _09259_ (.A0(_05389_),
    .A1(\tag_array.tag1[14][12] ),
    .S(_05592_),
    .X(_01013_));
 sky130_fd_sc_hd__mux2_1 _09260_ (.A0(_05391_),
    .A1(\tag_array.tag1[14][13] ),
    .S(_05592_),
    .X(_01014_));
 sky130_fd_sc_hd__mux2_1 _09261_ (.A0(_05393_),
    .A1(\tag_array.tag1[14][14] ),
    .S(_05592_),
    .X(_01015_));
 sky130_fd_sc_hd__mux2_1 _09262_ (.A0(_05395_),
    .A1(\tag_array.tag1[14][15] ),
    .S(_05592_),
    .X(_01016_));
 sky130_fd_sc_hd__mux2_1 _09263_ (.A0(_05397_),
    .A1(\tag_array.tag1[14][16] ),
    .S(_05592_),
    .X(_01017_));
 sky130_fd_sc_hd__mux2_1 _09264_ (.A0(_05399_),
    .A1(\tag_array.tag1[14][17] ),
    .S(_05592_),
    .X(_01018_));
 sky130_fd_sc_hd__mux2_1 _09265_ (.A0(_05401_),
    .A1(\tag_array.tag1[14][18] ),
    .S(_05592_),
    .X(_01019_));
 sky130_fd_sc_hd__mux2_1 _09266_ (.A0(_05403_),
    .A1(\tag_array.tag1[14][19] ),
    .S(_05592_),
    .X(_01020_));
 sky130_fd_sc_hd__mux2_1 _09267_ (.A0(_05405_),
    .A1(\tag_array.tag1[14][20] ),
    .S(_05592_),
    .X(_01021_));
 sky130_fd_sc_hd__mux2_1 _09268_ (.A0(_05407_),
    .A1(\tag_array.tag1[14][21] ),
    .S(_05592_),
    .X(_01022_));
 sky130_fd_sc_hd__mux2_1 _09269_ (.A0(_05409_),
    .A1(\tag_array.tag1[14][22] ),
    .S(_05592_),
    .X(_01023_));
 sky130_fd_sc_hd__mux2_1 _09270_ (.A0(_05411_),
    .A1(\tag_array.tag1[14][23] ),
    .S(_05592_),
    .X(_01024_));
 sky130_fd_sc_hd__mux2_1 _09271_ (.A0(_05413_),
    .A1(\tag_array.tag1[14][24] ),
    .S(_05592_),
    .X(_01025_));
 sky130_fd_sc_hd__mux2_1 _09272_ (.A0(_05365_),
    .A1(\tag_array.tag1[13][0] ),
    .S(_05593_),
    .X(_01026_));
 sky130_fd_sc_hd__mux2_1 _09273_ (.A0(_05367_),
    .A1(\tag_array.tag1[13][1] ),
    .S(_05593_),
    .X(_01027_));
 sky130_fd_sc_hd__mux2_1 _09274_ (.A0(_05369_),
    .A1(\tag_array.tag1[13][2] ),
    .S(_05593_),
    .X(_01028_));
 sky130_fd_sc_hd__mux2_1 _09275_ (.A0(_05371_),
    .A1(\tag_array.tag1[13][3] ),
    .S(_05593_),
    .X(_01029_));
 sky130_fd_sc_hd__mux2_1 _09276_ (.A0(_05373_),
    .A1(\tag_array.tag1[13][4] ),
    .S(_05593_),
    .X(_01030_));
 sky130_fd_sc_hd__mux2_1 _09277_ (.A0(_05375_),
    .A1(\tag_array.tag1[13][5] ),
    .S(_05593_),
    .X(_01031_));
 sky130_fd_sc_hd__mux2_1 _09278_ (.A0(_05377_),
    .A1(\tag_array.tag1[13][6] ),
    .S(_05593_),
    .X(_01032_));
 sky130_fd_sc_hd__mux2_1 _09279_ (.A0(_05379_),
    .A1(\tag_array.tag1[13][7] ),
    .S(_05593_),
    .X(_01033_));
 sky130_fd_sc_hd__mux2_1 _09280_ (.A0(_05381_),
    .A1(\tag_array.tag1[13][8] ),
    .S(_05593_),
    .X(_01034_));
 sky130_fd_sc_hd__mux2_1 _09281_ (.A0(_05383_),
    .A1(\tag_array.tag1[13][9] ),
    .S(_05593_),
    .X(_01035_));
 sky130_fd_sc_hd__mux2_1 _09282_ (.A0(_05385_),
    .A1(\tag_array.tag1[13][10] ),
    .S(_05593_),
    .X(_01036_));
 sky130_fd_sc_hd__mux2_1 _09283_ (.A0(_05387_),
    .A1(\tag_array.tag1[13][11] ),
    .S(_05593_),
    .X(_01037_));
 sky130_fd_sc_hd__mux2_1 _09284_ (.A0(_05389_),
    .A1(\tag_array.tag1[13][12] ),
    .S(_05593_),
    .X(_01038_));
 sky130_fd_sc_hd__mux2_1 _09285_ (.A0(_05391_),
    .A1(\tag_array.tag1[13][13] ),
    .S(_05593_),
    .X(_01039_));
 sky130_fd_sc_hd__mux2_1 _09286_ (.A0(_05393_),
    .A1(\tag_array.tag1[13][14] ),
    .S(_05593_),
    .X(_01040_));
 sky130_fd_sc_hd__mux2_1 _09287_ (.A0(_05395_),
    .A1(\tag_array.tag1[13][15] ),
    .S(_05593_),
    .X(_01041_));
 sky130_fd_sc_hd__mux2_1 _09288_ (.A0(_05397_),
    .A1(\tag_array.tag1[13][16] ),
    .S(_05593_),
    .X(_01042_));
 sky130_fd_sc_hd__mux2_1 _09289_ (.A0(_05399_),
    .A1(\tag_array.tag1[13][17] ),
    .S(_05593_),
    .X(_01043_));
 sky130_fd_sc_hd__mux2_1 _09290_ (.A0(_05401_),
    .A1(\tag_array.tag1[13][18] ),
    .S(_05593_),
    .X(_01044_));
 sky130_fd_sc_hd__mux2_1 _09291_ (.A0(_05403_),
    .A1(\tag_array.tag1[13][19] ),
    .S(_05593_),
    .X(_01045_));
 sky130_fd_sc_hd__mux2_1 _09292_ (.A0(_05405_),
    .A1(\tag_array.tag1[13][20] ),
    .S(_05593_),
    .X(_01046_));
 sky130_fd_sc_hd__mux2_1 _09293_ (.A0(_05407_),
    .A1(\tag_array.tag1[13][21] ),
    .S(_05593_),
    .X(_01047_));
 sky130_fd_sc_hd__mux2_1 _09294_ (.A0(_05409_),
    .A1(\tag_array.tag1[13][22] ),
    .S(_05593_),
    .X(_01048_));
 sky130_fd_sc_hd__mux2_1 _09295_ (.A0(_05411_),
    .A1(\tag_array.tag1[13][23] ),
    .S(_05593_),
    .X(_01049_));
 sky130_fd_sc_hd__mux2_1 _09296_ (.A0(_05413_),
    .A1(\tag_array.tag1[13][24] ),
    .S(_05593_),
    .X(_01050_));
 sky130_fd_sc_hd__mux2_1 _09297_ (.A0(_05365_),
    .A1(\tag_array.tag1[12][0] ),
    .S(_05594_),
    .X(_01051_));
 sky130_fd_sc_hd__mux2_1 _09298_ (.A0(_05367_),
    .A1(\tag_array.tag1[12][1] ),
    .S(_05594_),
    .X(_01052_));
 sky130_fd_sc_hd__mux2_1 _09299_ (.A0(_05369_),
    .A1(\tag_array.tag1[12][2] ),
    .S(_05594_),
    .X(_01053_));
 sky130_fd_sc_hd__mux2_1 _09300_ (.A0(_05371_),
    .A1(\tag_array.tag1[12][3] ),
    .S(_05594_),
    .X(_01054_));
 sky130_fd_sc_hd__mux2_1 _09301_ (.A0(_05373_),
    .A1(\tag_array.tag1[12][4] ),
    .S(_05594_),
    .X(_01055_));
 sky130_fd_sc_hd__mux2_1 _09302_ (.A0(_05375_),
    .A1(\tag_array.tag1[12][5] ),
    .S(_05594_),
    .X(_01056_));
 sky130_fd_sc_hd__mux2_1 _09303_ (.A0(_05377_),
    .A1(\tag_array.tag1[12][6] ),
    .S(_05594_),
    .X(_01057_));
 sky130_fd_sc_hd__mux2_1 _09304_ (.A0(_05379_),
    .A1(\tag_array.tag1[12][7] ),
    .S(_05594_),
    .X(_01058_));
 sky130_fd_sc_hd__mux2_1 _09305_ (.A0(_05381_),
    .A1(\tag_array.tag1[12][8] ),
    .S(_05594_),
    .X(_01059_));
 sky130_fd_sc_hd__mux2_1 _09306_ (.A0(_05383_),
    .A1(\tag_array.tag1[12][9] ),
    .S(_05594_),
    .X(_01060_));
 sky130_fd_sc_hd__mux2_1 _09307_ (.A0(_05385_),
    .A1(\tag_array.tag1[12][10] ),
    .S(_05594_),
    .X(_01061_));
 sky130_fd_sc_hd__mux2_1 _09308_ (.A0(_05387_),
    .A1(\tag_array.tag1[12][11] ),
    .S(_05594_),
    .X(_01062_));
 sky130_fd_sc_hd__mux2_1 _09309_ (.A0(_05389_),
    .A1(\tag_array.tag1[12][12] ),
    .S(_05594_),
    .X(_01063_));
 sky130_fd_sc_hd__mux2_1 _09310_ (.A0(_05391_),
    .A1(\tag_array.tag1[12][13] ),
    .S(_05594_),
    .X(_01064_));
 sky130_fd_sc_hd__mux2_1 _09311_ (.A0(_05393_),
    .A1(\tag_array.tag1[12][14] ),
    .S(_05594_),
    .X(_01065_));
 sky130_fd_sc_hd__mux2_1 _09312_ (.A0(_05395_),
    .A1(\tag_array.tag1[12][15] ),
    .S(_05594_),
    .X(_01066_));
 sky130_fd_sc_hd__mux2_1 _09313_ (.A0(_05397_),
    .A1(\tag_array.tag1[12][16] ),
    .S(_05594_),
    .X(_01067_));
 sky130_fd_sc_hd__mux2_1 _09314_ (.A0(_05399_),
    .A1(\tag_array.tag1[12][17] ),
    .S(_05594_),
    .X(_01068_));
 sky130_fd_sc_hd__mux2_1 _09315_ (.A0(_05401_),
    .A1(\tag_array.tag1[12][18] ),
    .S(_05594_),
    .X(_01069_));
 sky130_fd_sc_hd__mux2_1 _09316_ (.A0(_05403_),
    .A1(\tag_array.tag1[12][19] ),
    .S(_05594_),
    .X(_01070_));
 sky130_fd_sc_hd__mux2_1 _09317_ (.A0(_05405_),
    .A1(\tag_array.tag1[12][20] ),
    .S(_05594_),
    .X(_01071_));
 sky130_fd_sc_hd__mux2_1 _09318_ (.A0(_05407_),
    .A1(\tag_array.tag1[12][21] ),
    .S(_05594_),
    .X(_01072_));
 sky130_fd_sc_hd__mux2_1 _09319_ (.A0(_05409_),
    .A1(\tag_array.tag1[12][22] ),
    .S(_05594_),
    .X(_01073_));
 sky130_fd_sc_hd__mux2_1 _09320_ (.A0(_05411_),
    .A1(\tag_array.tag1[12][23] ),
    .S(_05594_),
    .X(_01074_));
 sky130_fd_sc_hd__mux2_1 _09321_ (.A0(_05413_),
    .A1(\tag_array.tag1[12][24] ),
    .S(_05594_),
    .X(_01075_));
 sky130_fd_sc_hd__or2_2 _09322_ (.A(_05414_),
    .B(_05552_),
    .X(_03123_));
 sky130_fd_sc_hd__mux2_1 _09323_ (.A0(_05420_),
    .A1(\data_array.data0[14][0] ),
    .S(_03123_),
    .X(_01076_));
 sky130_fd_sc_hd__mux2_1 _09324_ (.A0(_05422_),
    .A1(\data_array.data0[14][1] ),
    .S(_03123_),
    .X(_01077_));
 sky130_fd_sc_hd__mux2_1 _09325_ (.A0(_05424_),
    .A1(\data_array.data0[14][2] ),
    .S(_03123_),
    .X(_01078_));
 sky130_fd_sc_hd__mux2_1 _09326_ (.A0(_05426_),
    .A1(\data_array.data0[14][3] ),
    .S(_03123_),
    .X(_01079_));
 sky130_fd_sc_hd__mux2_1 _09327_ (.A0(_05428_),
    .A1(\data_array.data0[14][4] ),
    .S(_03123_),
    .X(_01080_));
 sky130_fd_sc_hd__mux2_1 _09328_ (.A0(_05430_),
    .A1(\data_array.data0[14][5] ),
    .S(_03123_),
    .X(_01081_));
 sky130_fd_sc_hd__mux2_1 _09329_ (.A0(_05432_),
    .A1(\data_array.data0[14][6] ),
    .S(_03123_),
    .X(_01082_));
 sky130_fd_sc_hd__mux2_1 _09330_ (.A0(_05434_),
    .A1(\data_array.data0[14][7] ),
    .S(_03123_),
    .X(_01083_));
 sky130_fd_sc_hd__mux2_1 _09331_ (.A0(_05436_),
    .A1(\data_array.data0[14][8] ),
    .S(_03123_),
    .X(_01084_));
 sky130_fd_sc_hd__mux2_1 _09332_ (.A0(_05438_),
    .A1(\data_array.data0[14][9] ),
    .S(_03123_),
    .X(_01085_));
 sky130_fd_sc_hd__mux2_1 _09333_ (.A0(_05440_),
    .A1(\data_array.data0[14][10] ),
    .S(_03123_),
    .X(_01086_));
 sky130_fd_sc_hd__mux2_1 _09334_ (.A0(_05442_),
    .A1(\data_array.data0[14][11] ),
    .S(_03123_),
    .X(_01087_));
 sky130_fd_sc_hd__mux2_1 _09335_ (.A0(_05444_),
    .A1(\data_array.data0[14][12] ),
    .S(_03123_),
    .X(_01088_));
 sky130_fd_sc_hd__mux2_1 _09336_ (.A0(_05446_),
    .A1(\data_array.data0[14][13] ),
    .S(_03123_),
    .X(_01089_));
 sky130_fd_sc_hd__mux2_1 _09337_ (.A0(_05448_),
    .A1(\data_array.data0[14][14] ),
    .S(_03123_),
    .X(_01090_));
 sky130_fd_sc_hd__mux2_1 _09338_ (.A0(_05450_),
    .A1(\data_array.data0[14][15] ),
    .S(_03123_),
    .X(_01091_));
 sky130_fd_sc_hd__mux2_1 _09339_ (.A0(_05452_),
    .A1(\data_array.data0[14][16] ),
    .S(_03123_),
    .X(_01092_));
 sky130_fd_sc_hd__mux2_1 _09340_ (.A0(_05454_),
    .A1(\data_array.data0[14][17] ),
    .S(_03123_),
    .X(_01093_));
 sky130_fd_sc_hd__mux2_1 _09341_ (.A0(_05456_),
    .A1(\data_array.data0[14][18] ),
    .S(_03123_),
    .X(_01094_));
 sky130_fd_sc_hd__mux2_1 _09342_ (.A0(_05458_),
    .A1(\data_array.data0[14][19] ),
    .S(_03123_),
    .X(_01095_));
 sky130_fd_sc_hd__mux2_1 _09343_ (.A0(_05460_),
    .A1(\data_array.data0[14][20] ),
    .S(_03123_),
    .X(_01096_));
 sky130_fd_sc_hd__mux2_1 _09344_ (.A0(_05462_),
    .A1(\data_array.data0[14][21] ),
    .S(_03123_),
    .X(_01097_));
 sky130_fd_sc_hd__mux2_1 _09345_ (.A0(_05464_),
    .A1(\data_array.data0[14][22] ),
    .S(_03123_),
    .X(_01098_));
 sky130_fd_sc_hd__mux2_1 _09346_ (.A0(_05466_),
    .A1(\data_array.data0[14][23] ),
    .S(_03123_),
    .X(_01099_));
 sky130_fd_sc_hd__mux2_1 _09347_ (.A0(_05468_),
    .A1(\data_array.data0[14][24] ),
    .S(_03123_),
    .X(_01100_));
 sky130_fd_sc_hd__mux2_1 _09348_ (.A0(_05470_),
    .A1(\data_array.data0[14][25] ),
    .S(_03123_),
    .X(_01101_));
 sky130_fd_sc_hd__mux2_1 _09349_ (.A0(_05472_),
    .A1(\data_array.data0[14][26] ),
    .S(_03123_),
    .X(_01102_));
 sky130_fd_sc_hd__mux2_1 _09350_ (.A0(_05474_),
    .A1(\data_array.data0[14][27] ),
    .S(_03123_),
    .X(_01103_));
 sky130_fd_sc_hd__mux2_1 _09351_ (.A0(_05476_),
    .A1(\data_array.data0[14][28] ),
    .S(_03123_),
    .X(_01104_));
 sky130_fd_sc_hd__mux2_1 _09352_ (.A0(_05478_),
    .A1(\data_array.data0[14][29] ),
    .S(_03123_),
    .X(_01105_));
 sky130_fd_sc_hd__mux2_1 _09353_ (.A0(_05480_),
    .A1(\data_array.data0[14][30] ),
    .S(_03123_),
    .X(_01106_));
 sky130_fd_sc_hd__mux2_1 _09354_ (.A0(_05482_),
    .A1(\data_array.data0[14][31] ),
    .S(_03123_),
    .X(_01107_));
 sky130_fd_sc_hd__mux2_1 _09355_ (.A0(_05484_),
    .A1(\data_array.data0[14][32] ),
    .S(_03123_),
    .X(_01108_));
 sky130_fd_sc_hd__mux2_1 _09356_ (.A0(_05486_),
    .A1(\data_array.data0[14][33] ),
    .S(_03123_),
    .X(_01109_));
 sky130_fd_sc_hd__mux2_1 _09357_ (.A0(_05488_),
    .A1(\data_array.data0[14][34] ),
    .S(_03123_),
    .X(_01110_));
 sky130_fd_sc_hd__mux2_1 _09358_ (.A0(_05490_),
    .A1(\data_array.data0[14][35] ),
    .S(_03123_),
    .X(_01111_));
 sky130_fd_sc_hd__mux2_1 _09359_ (.A0(_05492_),
    .A1(\data_array.data0[14][36] ),
    .S(_03123_),
    .X(_01112_));
 sky130_fd_sc_hd__mux2_1 _09360_ (.A0(_05494_),
    .A1(\data_array.data0[14][37] ),
    .S(_03123_),
    .X(_01113_));
 sky130_fd_sc_hd__mux2_1 _09361_ (.A0(_05496_),
    .A1(\data_array.data0[14][38] ),
    .S(_03123_),
    .X(_01114_));
 sky130_fd_sc_hd__mux2_1 _09362_ (.A0(_05498_),
    .A1(\data_array.data0[14][39] ),
    .S(_03123_),
    .X(_01115_));
 sky130_fd_sc_hd__mux2_1 _09363_ (.A0(_05500_),
    .A1(\data_array.data0[14][40] ),
    .S(_03123_),
    .X(_01116_));
 sky130_fd_sc_hd__mux2_1 _09364_ (.A0(_05502_),
    .A1(\data_array.data0[14][41] ),
    .S(_03123_),
    .X(_01117_));
 sky130_fd_sc_hd__mux2_1 _09365_ (.A0(_05504_),
    .A1(\data_array.data0[14][42] ),
    .S(_03123_),
    .X(_01118_));
 sky130_fd_sc_hd__mux2_1 _09366_ (.A0(_05506_),
    .A1(\data_array.data0[14][43] ),
    .S(_03123_),
    .X(_01119_));
 sky130_fd_sc_hd__mux2_1 _09367_ (.A0(_05508_),
    .A1(\data_array.data0[14][44] ),
    .S(_03123_),
    .X(_01120_));
 sky130_fd_sc_hd__mux2_1 _09368_ (.A0(_05510_),
    .A1(\data_array.data0[14][45] ),
    .S(_03123_),
    .X(_01121_));
 sky130_fd_sc_hd__mux2_1 _09369_ (.A0(_05512_),
    .A1(\data_array.data0[14][46] ),
    .S(_03123_),
    .X(_01122_));
 sky130_fd_sc_hd__mux2_1 _09370_ (.A0(_05514_),
    .A1(\data_array.data0[14][47] ),
    .S(_03123_),
    .X(_01123_));
 sky130_fd_sc_hd__mux2_1 _09371_ (.A0(_05516_),
    .A1(\data_array.data0[14][48] ),
    .S(_03123_),
    .X(_01124_));
 sky130_fd_sc_hd__mux2_1 _09372_ (.A0(_05518_),
    .A1(\data_array.data0[14][49] ),
    .S(_03123_),
    .X(_01125_));
 sky130_fd_sc_hd__mux2_1 _09373_ (.A0(_05520_),
    .A1(\data_array.data0[14][50] ),
    .S(_03123_),
    .X(_01126_));
 sky130_fd_sc_hd__mux2_1 _09374_ (.A0(_05522_),
    .A1(\data_array.data0[14][51] ),
    .S(_03123_),
    .X(_01127_));
 sky130_fd_sc_hd__mux2_1 _09375_ (.A0(_05524_),
    .A1(\data_array.data0[14][52] ),
    .S(_03123_),
    .X(_01128_));
 sky130_fd_sc_hd__mux2_1 _09376_ (.A0(_05526_),
    .A1(\data_array.data0[14][53] ),
    .S(_03123_),
    .X(_01129_));
 sky130_fd_sc_hd__mux2_1 _09377_ (.A0(_05528_),
    .A1(\data_array.data0[14][54] ),
    .S(_03123_),
    .X(_01130_));
 sky130_fd_sc_hd__mux2_1 _09378_ (.A0(_05530_),
    .A1(\data_array.data0[14][55] ),
    .S(_03123_),
    .X(_01131_));
 sky130_fd_sc_hd__mux2_1 _09379_ (.A0(_05532_),
    .A1(\data_array.data0[14][56] ),
    .S(_03123_),
    .X(_01132_));
 sky130_fd_sc_hd__mux2_1 _09380_ (.A0(_05534_),
    .A1(\data_array.data0[14][57] ),
    .S(_03123_),
    .X(_01133_));
 sky130_fd_sc_hd__mux2_1 _09381_ (.A0(_05536_),
    .A1(\data_array.data0[14][58] ),
    .S(_03123_),
    .X(_01134_));
 sky130_fd_sc_hd__mux2_1 _09382_ (.A0(_05538_),
    .A1(\data_array.data0[14][59] ),
    .S(_03123_),
    .X(_01135_));
 sky130_fd_sc_hd__mux2_1 _09383_ (.A0(_05540_),
    .A1(\data_array.data0[14][60] ),
    .S(_03123_),
    .X(_01136_));
 sky130_fd_sc_hd__mux2_1 _09384_ (.A0(_05542_),
    .A1(\data_array.data0[14][61] ),
    .S(_03123_),
    .X(_01137_));
 sky130_fd_sc_hd__mux2_1 _09385_ (.A0(_05544_),
    .A1(\data_array.data0[14][62] ),
    .S(_03123_),
    .X(_01138_));
 sky130_fd_sc_hd__mux2_1 _09386_ (.A0(_05546_),
    .A1(\data_array.data0[14][63] ),
    .S(_03123_),
    .X(_01139_));
 sky130_fd_sc_hd__mux2_1 _09387_ (.A0(_05356_),
    .A1(\lru_array.lru_mem[6] ),
    .S(_05575_),
    .X(_01140_));
 sky130_fd_sc_hd__mux2_1 _09388_ (.A0(_05356_),
    .A1(\lru_array.lru_mem[7] ),
    .S(_05572_),
    .X(_01141_));
 sky130_fd_sc_hd__mux2_1 _09389_ (.A0(_05420_),
    .A1(\data_array.data1[9][0] ),
    .S(_05591_),
    .X(_01142_));
 sky130_fd_sc_hd__mux2_1 _09390_ (.A0(_05422_),
    .A1(\data_array.data1[9][1] ),
    .S(_05591_),
    .X(_01143_));
 sky130_fd_sc_hd__mux2_1 _09391_ (.A0(_05424_),
    .A1(\data_array.data1[9][2] ),
    .S(_05591_),
    .X(_01144_));
 sky130_fd_sc_hd__mux2_1 _09392_ (.A0(_05426_),
    .A1(\data_array.data1[9][3] ),
    .S(_05591_),
    .X(_01145_));
 sky130_fd_sc_hd__mux2_1 _09393_ (.A0(_05428_),
    .A1(\data_array.data1[9][4] ),
    .S(_05591_),
    .X(_01146_));
 sky130_fd_sc_hd__mux2_1 _09394_ (.A0(_05430_),
    .A1(\data_array.data1[9][5] ),
    .S(_05591_),
    .X(_01147_));
 sky130_fd_sc_hd__mux2_1 _09395_ (.A0(_05432_),
    .A1(\data_array.data1[9][6] ),
    .S(_05591_),
    .X(_01148_));
 sky130_fd_sc_hd__mux2_1 _09396_ (.A0(_05434_),
    .A1(\data_array.data1[9][7] ),
    .S(_05591_),
    .X(_01149_));
 sky130_fd_sc_hd__mux2_1 _09397_ (.A0(_05436_),
    .A1(\data_array.data1[9][8] ),
    .S(_05591_),
    .X(_01150_));
 sky130_fd_sc_hd__mux2_1 _09398_ (.A0(_05438_),
    .A1(\data_array.data1[9][9] ),
    .S(_05591_),
    .X(_01151_));
 sky130_fd_sc_hd__mux2_1 _09399_ (.A0(_05440_),
    .A1(\data_array.data1[9][10] ),
    .S(_05591_),
    .X(_01152_));
 sky130_fd_sc_hd__mux2_1 _09400_ (.A0(_05442_),
    .A1(\data_array.data1[9][11] ),
    .S(_05591_),
    .X(_01153_));
 sky130_fd_sc_hd__mux2_1 _09401_ (.A0(_05444_),
    .A1(\data_array.data1[9][12] ),
    .S(_05591_),
    .X(_01154_));
 sky130_fd_sc_hd__mux2_1 _09402_ (.A0(_05446_),
    .A1(\data_array.data1[9][13] ),
    .S(_05591_),
    .X(_01155_));
 sky130_fd_sc_hd__mux2_1 _09403_ (.A0(_05448_),
    .A1(\data_array.data1[9][14] ),
    .S(_05591_),
    .X(_01156_));
 sky130_fd_sc_hd__mux2_1 _09404_ (.A0(_05450_),
    .A1(\data_array.data1[9][15] ),
    .S(_05591_),
    .X(_01157_));
 sky130_fd_sc_hd__mux2_1 _09405_ (.A0(_05452_),
    .A1(\data_array.data1[9][16] ),
    .S(_05591_),
    .X(_01158_));
 sky130_fd_sc_hd__mux2_1 _09406_ (.A0(_05454_),
    .A1(\data_array.data1[9][17] ),
    .S(_05591_),
    .X(_01159_));
 sky130_fd_sc_hd__mux2_1 _09407_ (.A0(_05456_),
    .A1(\data_array.data1[9][18] ),
    .S(_05591_),
    .X(_01160_));
 sky130_fd_sc_hd__mux2_1 _09408_ (.A0(_05458_),
    .A1(\data_array.data1[9][19] ),
    .S(_05591_),
    .X(_01161_));
 sky130_fd_sc_hd__mux2_1 _09409_ (.A0(_05460_),
    .A1(\data_array.data1[9][20] ),
    .S(_05591_),
    .X(_01162_));
 sky130_fd_sc_hd__mux2_1 _09410_ (.A0(_05462_),
    .A1(\data_array.data1[9][21] ),
    .S(_05591_),
    .X(_01163_));
 sky130_fd_sc_hd__mux2_1 _09411_ (.A0(_05464_),
    .A1(\data_array.data1[9][22] ),
    .S(_05591_),
    .X(_01164_));
 sky130_fd_sc_hd__mux2_1 _09412_ (.A0(_05466_),
    .A1(\data_array.data1[9][23] ),
    .S(_05591_),
    .X(_01165_));
 sky130_fd_sc_hd__mux2_1 _09413_ (.A0(_05468_),
    .A1(\data_array.data1[9][24] ),
    .S(_05591_),
    .X(_01166_));
 sky130_fd_sc_hd__mux2_1 _09414_ (.A0(_05470_),
    .A1(\data_array.data1[9][25] ),
    .S(_05591_),
    .X(_01167_));
 sky130_fd_sc_hd__mux2_1 _09415_ (.A0(_05472_),
    .A1(\data_array.data1[9][26] ),
    .S(_05591_),
    .X(_01168_));
 sky130_fd_sc_hd__mux2_1 _09416_ (.A0(_05474_),
    .A1(\data_array.data1[9][27] ),
    .S(_05591_),
    .X(_01169_));
 sky130_fd_sc_hd__mux2_1 _09417_ (.A0(_05476_),
    .A1(\data_array.data1[9][28] ),
    .S(_05591_),
    .X(_01170_));
 sky130_fd_sc_hd__mux2_1 _09418_ (.A0(_05478_),
    .A1(\data_array.data1[9][29] ),
    .S(_05591_),
    .X(_01171_));
 sky130_fd_sc_hd__mux2_1 _09419_ (.A0(_05480_),
    .A1(\data_array.data1[9][30] ),
    .S(_05591_),
    .X(_01172_));
 sky130_fd_sc_hd__mux2_1 _09420_ (.A0(_05482_),
    .A1(\data_array.data1[9][31] ),
    .S(_05591_),
    .X(_01173_));
 sky130_fd_sc_hd__mux2_1 _09421_ (.A0(_05484_),
    .A1(\data_array.data1[9][32] ),
    .S(_05591_),
    .X(_01174_));
 sky130_fd_sc_hd__mux2_1 _09422_ (.A0(_05486_),
    .A1(\data_array.data1[9][33] ),
    .S(_05591_),
    .X(_01175_));
 sky130_fd_sc_hd__mux2_1 _09423_ (.A0(_05488_),
    .A1(\data_array.data1[9][34] ),
    .S(_05591_),
    .X(_01176_));
 sky130_fd_sc_hd__mux2_1 _09424_ (.A0(_05490_),
    .A1(\data_array.data1[9][35] ),
    .S(_05591_),
    .X(_01177_));
 sky130_fd_sc_hd__mux2_1 _09425_ (.A0(_05492_),
    .A1(\data_array.data1[9][36] ),
    .S(_05591_),
    .X(_01178_));
 sky130_fd_sc_hd__mux2_1 _09426_ (.A0(_05494_),
    .A1(\data_array.data1[9][37] ),
    .S(_05591_),
    .X(_01179_));
 sky130_fd_sc_hd__mux2_1 _09427_ (.A0(_05496_),
    .A1(\data_array.data1[9][38] ),
    .S(_05591_),
    .X(_01180_));
 sky130_fd_sc_hd__mux2_1 _09428_ (.A0(_05498_),
    .A1(\data_array.data1[9][39] ),
    .S(_05591_),
    .X(_01181_));
 sky130_fd_sc_hd__mux2_1 _09429_ (.A0(_05500_),
    .A1(\data_array.data1[9][40] ),
    .S(_05591_),
    .X(_01182_));
 sky130_fd_sc_hd__mux2_1 _09430_ (.A0(_05502_),
    .A1(\data_array.data1[9][41] ),
    .S(_05591_),
    .X(_01183_));
 sky130_fd_sc_hd__mux2_1 _09431_ (.A0(_05504_),
    .A1(\data_array.data1[9][42] ),
    .S(_05591_),
    .X(_01184_));
 sky130_fd_sc_hd__mux2_1 _09432_ (.A0(_05506_),
    .A1(\data_array.data1[9][43] ),
    .S(_05591_),
    .X(_01185_));
 sky130_fd_sc_hd__mux2_1 _09433_ (.A0(_05508_),
    .A1(\data_array.data1[9][44] ),
    .S(_05591_),
    .X(_01186_));
 sky130_fd_sc_hd__mux2_1 _09434_ (.A0(_05510_),
    .A1(\data_array.data1[9][45] ),
    .S(_05591_),
    .X(_01187_));
 sky130_fd_sc_hd__mux2_1 _09435_ (.A0(_05512_),
    .A1(\data_array.data1[9][46] ),
    .S(_05591_),
    .X(_01188_));
 sky130_fd_sc_hd__mux2_1 _09436_ (.A0(_05514_),
    .A1(\data_array.data1[9][47] ),
    .S(_05591_),
    .X(_01189_));
 sky130_fd_sc_hd__mux2_1 _09437_ (.A0(_05516_),
    .A1(\data_array.data1[9][48] ),
    .S(_05591_),
    .X(_01190_));
 sky130_fd_sc_hd__mux2_1 _09438_ (.A0(_05518_),
    .A1(\data_array.data1[9][49] ),
    .S(_05591_),
    .X(_01191_));
 sky130_fd_sc_hd__mux2_1 _09439_ (.A0(_05520_),
    .A1(\data_array.data1[9][50] ),
    .S(_05591_),
    .X(_01192_));
 sky130_fd_sc_hd__mux2_1 _09440_ (.A0(_05522_),
    .A1(\data_array.data1[9][51] ),
    .S(_05591_),
    .X(_01193_));
 sky130_fd_sc_hd__mux2_1 _09441_ (.A0(_05524_),
    .A1(\data_array.data1[9][52] ),
    .S(_05591_),
    .X(_01194_));
 sky130_fd_sc_hd__mux2_1 _09442_ (.A0(_05526_),
    .A1(\data_array.data1[9][53] ),
    .S(_05591_),
    .X(_01195_));
 sky130_fd_sc_hd__mux2_1 _09443_ (.A0(_05528_),
    .A1(\data_array.data1[9][54] ),
    .S(_05591_),
    .X(_01196_));
 sky130_fd_sc_hd__mux2_1 _09444_ (.A0(_05530_),
    .A1(\data_array.data1[9][55] ),
    .S(_05591_),
    .X(_01197_));
 sky130_fd_sc_hd__mux2_1 _09445_ (.A0(_05532_),
    .A1(\data_array.data1[9][56] ),
    .S(_05591_),
    .X(_01198_));
 sky130_fd_sc_hd__mux2_1 _09446_ (.A0(_05534_),
    .A1(\data_array.data1[9][57] ),
    .S(_05591_),
    .X(_01199_));
 sky130_fd_sc_hd__mux2_1 _09447_ (.A0(_05536_),
    .A1(\data_array.data1[9][58] ),
    .S(_05591_),
    .X(_01200_));
 sky130_fd_sc_hd__mux2_1 _09448_ (.A0(_05538_),
    .A1(\data_array.data1[9][59] ),
    .S(_05591_),
    .X(_01201_));
 sky130_fd_sc_hd__mux2_1 _09449_ (.A0(_05540_),
    .A1(\data_array.data1[9][60] ),
    .S(_05591_),
    .X(_01202_));
 sky130_fd_sc_hd__mux2_1 _09450_ (.A0(_05542_),
    .A1(\data_array.data1[9][61] ),
    .S(_05591_),
    .X(_01203_));
 sky130_fd_sc_hd__mux2_1 _09451_ (.A0(_05544_),
    .A1(\data_array.data1[9][62] ),
    .S(_05591_),
    .X(_01204_));
 sky130_fd_sc_hd__mux2_1 _09452_ (.A0(_05546_),
    .A1(\data_array.data1[9][63] ),
    .S(_05591_),
    .X(_01205_));
 sky130_fd_sc_hd__mux2_1 _09453_ (.A0(_05356_),
    .A1(\lru_array.lru_mem[8] ),
    .S(_05570_),
    .X(_01206_));
 sky130_fd_sc_hd__mux2_1 _09454_ (.A0(_05356_),
    .A1(\lru_array.lru_mem[0] ),
    .S(_05568_),
    .X(_01207_));
 sky130_fd_sc_hd__mux2_1 _09455_ (.A0(_05356_),
    .A1(\lru_array.lru_mem[15] ),
    .S(_05596_),
    .X(_01208_));
 sky130_fd_sc_hd__mux2_1 _09456_ (.A0(_05356_),
    .A1(\lru_array.lru_mem[10] ),
    .S(_05566_),
    .X(_01209_));
 sky130_fd_sc_hd__mux2_1 _09457_ (.A0(_05356_),
    .A1(\lru_array.lru_mem[1] ),
    .S(_05588_),
    .X(_01210_));
 sky130_fd_sc_hd__mux2_1 _09458_ (.A0(_05356_),
    .A1(\lru_array.lru_mem[11] ),
    .S(_05564_),
    .X(_01211_));
 sky130_fd_sc_hd__mux2_1 _09459_ (.A0(_05365_),
    .A1(\tag_array.tag1[11][0] ),
    .S(_05551_),
    .X(_01212_));
 sky130_fd_sc_hd__mux2_1 _09460_ (.A0(_05367_),
    .A1(\tag_array.tag1[11][1] ),
    .S(_05551_),
    .X(_01213_));
 sky130_fd_sc_hd__mux2_1 _09461_ (.A0(_05369_),
    .A1(\tag_array.tag1[11][2] ),
    .S(_05551_),
    .X(_01214_));
 sky130_fd_sc_hd__mux2_1 _09462_ (.A0(_05371_),
    .A1(\tag_array.tag1[11][3] ),
    .S(_05551_),
    .X(_01215_));
 sky130_fd_sc_hd__mux2_1 _09463_ (.A0(_05373_),
    .A1(\tag_array.tag1[11][4] ),
    .S(_05551_),
    .X(_01216_));
 sky130_fd_sc_hd__mux2_1 _09464_ (.A0(_05375_),
    .A1(\tag_array.tag1[11][5] ),
    .S(_05551_),
    .X(_01217_));
 sky130_fd_sc_hd__mux2_1 _09465_ (.A0(_05377_),
    .A1(\tag_array.tag1[11][6] ),
    .S(_05551_),
    .X(_01218_));
 sky130_fd_sc_hd__mux2_1 _09466_ (.A0(_05379_),
    .A1(\tag_array.tag1[11][7] ),
    .S(_05551_),
    .X(_01219_));
 sky130_fd_sc_hd__mux2_1 _09467_ (.A0(_05381_),
    .A1(\tag_array.tag1[11][8] ),
    .S(_05551_),
    .X(_01220_));
 sky130_fd_sc_hd__mux2_1 _09468_ (.A0(_05383_),
    .A1(\tag_array.tag1[11][9] ),
    .S(_05551_),
    .X(_01221_));
 sky130_fd_sc_hd__mux2_1 _09469_ (.A0(_05385_),
    .A1(\tag_array.tag1[11][10] ),
    .S(_05551_),
    .X(_01222_));
 sky130_fd_sc_hd__mux2_1 _09470_ (.A0(_05387_),
    .A1(\tag_array.tag1[11][11] ),
    .S(_05551_),
    .X(_01223_));
 sky130_fd_sc_hd__mux2_1 _09471_ (.A0(_05389_),
    .A1(\tag_array.tag1[11][12] ),
    .S(_05551_),
    .X(_01224_));
 sky130_fd_sc_hd__mux2_1 _09472_ (.A0(_05391_),
    .A1(\tag_array.tag1[11][13] ),
    .S(_05551_),
    .X(_01225_));
 sky130_fd_sc_hd__mux2_1 _09473_ (.A0(_05393_),
    .A1(\tag_array.tag1[11][14] ),
    .S(_05551_),
    .X(_01226_));
 sky130_fd_sc_hd__mux2_1 _09474_ (.A0(_05395_),
    .A1(\tag_array.tag1[11][15] ),
    .S(_05551_),
    .X(_01227_));
 sky130_fd_sc_hd__mux2_1 _09475_ (.A0(_05397_),
    .A1(\tag_array.tag1[11][16] ),
    .S(_05551_),
    .X(_01228_));
 sky130_fd_sc_hd__mux2_1 _09476_ (.A0(_05399_),
    .A1(\tag_array.tag1[11][17] ),
    .S(_05551_),
    .X(_01229_));
 sky130_fd_sc_hd__mux2_1 _09477_ (.A0(_05401_),
    .A1(\tag_array.tag1[11][18] ),
    .S(_05551_),
    .X(_01230_));
 sky130_fd_sc_hd__mux2_1 _09478_ (.A0(_05403_),
    .A1(\tag_array.tag1[11][19] ),
    .S(_05551_),
    .X(_01231_));
 sky130_fd_sc_hd__mux2_1 _09479_ (.A0(_05405_),
    .A1(\tag_array.tag1[11][20] ),
    .S(_05551_),
    .X(_01232_));
 sky130_fd_sc_hd__mux2_1 _09480_ (.A0(_05407_),
    .A1(\tag_array.tag1[11][21] ),
    .S(_05551_),
    .X(_01233_));
 sky130_fd_sc_hd__mux2_1 _09481_ (.A0(_05409_),
    .A1(\tag_array.tag1[11][22] ),
    .S(_05551_),
    .X(_01234_));
 sky130_fd_sc_hd__mux2_1 _09482_ (.A0(_05411_),
    .A1(\tag_array.tag1[11][23] ),
    .S(_05551_),
    .X(_01235_));
 sky130_fd_sc_hd__mux2_1 _09483_ (.A0(_05413_),
    .A1(\tag_array.tag1[11][24] ),
    .S(_05551_),
    .X(_01236_));
 sky130_fd_sc_hd__mux2_1 _09484_ (.A0(_05365_),
    .A1(\tag_array.tag0[11][0] ),
    .S(_05565_),
    .X(_01237_));
 sky130_fd_sc_hd__mux2_1 _09485_ (.A0(_05367_),
    .A1(\tag_array.tag0[11][1] ),
    .S(_05565_),
    .X(_01238_));
 sky130_fd_sc_hd__mux2_1 _09486_ (.A0(_05369_),
    .A1(\tag_array.tag0[11][2] ),
    .S(_05565_),
    .X(_01239_));
 sky130_fd_sc_hd__mux2_1 _09487_ (.A0(_05371_),
    .A1(\tag_array.tag0[11][3] ),
    .S(_05565_),
    .X(_01240_));
 sky130_fd_sc_hd__mux2_1 _09488_ (.A0(_05373_),
    .A1(\tag_array.tag0[11][4] ),
    .S(_05565_),
    .X(_01241_));
 sky130_fd_sc_hd__mux2_1 _09489_ (.A0(_05375_),
    .A1(\tag_array.tag0[11][5] ),
    .S(_05565_),
    .X(_01242_));
 sky130_fd_sc_hd__mux2_1 _09490_ (.A0(_05377_),
    .A1(\tag_array.tag0[11][6] ),
    .S(_05565_),
    .X(_01243_));
 sky130_fd_sc_hd__mux2_1 _09491_ (.A0(_05379_),
    .A1(\tag_array.tag0[11][7] ),
    .S(_05565_),
    .X(_01244_));
 sky130_fd_sc_hd__mux2_1 _09492_ (.A0(_05381_),
    .A1(\tag_array.tag0[11][8] ),
    .S(_05565_),
    .X(_01245_));
 sky130_fd_sc_hd__mux2_1 _09493_ (.A0(_05383_),
    .A1(\tag_array.tag0[11][9] ),
    .S(_05565_),
    .X(_01246_));
 sky130_fd_sc_hd__mux2_1 _09494_ (.A0(_05385_),
    .A1(\tag_array.tag0[11][10] ),
    .S(_05565_),
    .X(_01247_));
 sky130_fd_sc_hd__mux2_1 _09495_ (.A0(_05387_),
    .A1(\tag_array.tag0[11][11] ),
    .S(_05565_),
    .X(_01248_));
 sky130_fd_sc_hd__mux2_1 _09496_ (.A0(_05389_),
    .A1(\tag_array.tag0[11][12] ),
    .S(_05565_),
    .X(_01249_));
 sky130_fd_sc_hd__mux2_1 _09497_ (.A0(_05391_),
    .A1(\tag_array.tag0[11][13] ),
    .S(_05565_),
    .X(_01250_));
 sky130_fd_sc_hd__mux2_1 _09498_ (.A0(_05393_),
    .A1(\tag_array.tag0[11][14] ),
    .S(_05565_),
    .X(_01251_));
 sky130_fd_sc_hd__mux2_1 _09499_ (.A0(_05395_),
    .A1(\tag_array.tag0[11][15] ),
    .S(_05565_),
    .X(_01252_));
 sky130_fd_sc_hd__mux2_1 _09500_ (.A0(_05397_),
    .A1(\tag_array.tag0[11][16] ),
    .S(_05565_),
    .X(_01253_));
 sky130_fd_sc_hd__mux2_1 _09501_ (.A0(_05399_),
    .A1(\tag_array.tag0[11][17] ),
    .S(_05565_),
    .X(_01254_));
 sky130_fd_sc_hd__mux2_1 _09502_ (.A0(_05401_),
    .A1(\tag_array.tag0[11][18] ),
    .S(_05565_),
    .X(_01255_));
 sky130_fd_sc_hd__mux2_1 _09503_ (.A0(_05403_),
    .A1(\tag_array.tag0[11][19] ),
    .S(_05565_),
    .X(_01256_));
 sky130_fd_sc_hd__mux2_1 _09504_ (.A0(_05405_),
    .A1(\tag_array.tag0[11][20] ),
    .S(_05565_),
    .X(_01257_));
 sky130_fd_sc_hd__mux2_1 _09505_ (.A0(_05407_),
    .A1(\tag_array.tag0[11][21] ),
    .S(_05565_),
    .X(_01258_));
 sky130_fd_sc_hd__mux2_1 _09506_ (.A0(_05409_),
    .A1(\tag_array.tag0[11][22] ),
    .S(_05565_),
    .X(_01259_));
 sky130_fd_sc_hd__mux2_1 _09507_ (.A0(_05411_),
    .A1(\tag_array.tag0[11][23] ),
    .S(_05565_),
    .X(_01260_));
 sky130_fd_sc_hd__mux2_1 _09508_ (.A0(_05413_),
    .A1(\tag_array.tag0[11][24] ),
    .S(_05565_),
    .X(_01261_));
 sky130_fd_sc_hd__mux2_1 _09509_ (.A0(_05365_),
    .A1(\tag_array.tag0[10][0] ),
    .S(_05567_),
    .X(_01262_));
 sky130_fd_sc_hd__mux2_1 _09510_ (.A0(_05367_),
    .A1(\tag_array.tag0[10][1] ),
    .S(_05567_),
    .X(_01263_));
 sky130_fd_sc_hd__mux2_1 _09511_ (.A0(_05369_),
    .A1(\tag_array.tag0[10][2] ),
    .S(_05567_),
    .X(_01264_));
 sky130_fd_sc_hd__mux2_1 _09512_ (.A0(_05371_),
    .A1(\tag_array.tag0[10][3] ),
    .S(_05567_),
    .X(_01265_));
 sky130_fd_sc_hd__mux2_1 _09513_ (.A0(_05373_),
    .A1(\tag_array.tag0[10][4] ),
    .S(_05567_),
    .X(_01266_));
 sky130_fd_sc_hd__mux2_1 _09514_ (.A0(_05375_),
    .A1(\tag_array.tag0[10][5] ),
    .S(_05567_),
    .X(_01267_));
 sky130_fd_sc_hd__mux2_1 _09515_ (.A0(_05377_),
    .A1(\tag_array.tag0[10][6] ),
    .S(_05567_),
    .X(_01268_));
 sky130_fd_sc_hd__mux2_1 _09516_ (.A0(_05379_),
    .A1(\tag_array.tag0[10][7] ),
    .S(_05567_),
    .X(_01269_));
 sky130_fd_sc_hd__mux2_1 _09517_ (.A0(_05381_),
    .A1(\tag_array.tag0[10][8] ),
    .S(_05567_),
    .X(_01270_));
 sky130_fd_sc_hd__mux2_1 _09518_ (.A0(_05383_),
    .A1(\tag_array.tag0[10][9] ),
    .S(_05567_),
    .X(_01271_));
 sky130_fd_sc_hd__mux2_1 _09519_ (.A0(_05385_),
    .A1(\tag_array.tag0[10][10] ),
    .S(_05567_),
    .X(_01272_));
 sky130_fd_sc_hd__mux2_1 _09520_ (.A0(_05387_),
    .A1(\tag_array.tag0[10][11] ),
    .S(_05567_),
    .X(_01273_));
 sky130_fd_sc_hd__mux2_1 _09521_ (.A0(_05389_),
    .A1(\tag_array.tag0[10][12] ),
    .S(_05567_),
    .X(_01274_));
 sky130_fd_sc_hd__mux2_1 _09522_ (.A0(_05391_),
    .A1(\tag_array.tag0[10][13] ),
    .S(_05567_),
    .X(_01275_));
 sky130_fd_sc_hd__mux2_1 _09523_ (.A0(_05393_),
    .A1(\tag_array.tag0[10][14] ),
    .S(_05567_),
    .X(_01276_));
 sky130_fd_sc_hd__mux2_1 _09524_ (.A0(_05395_),
    .A1(\tag_array.tag0[10][15] ),
    .S(_05567_),
    .X(_01277_));
 sky130_fd_sc_hd__mux2_1 _09525_ (.A0(_05397_),
    .A1(\tag_array.tag0[10][16] ),
    .S(_05567_),
    .X(_01278_));
 sky130_fd_sc_hd__mux2_1 _09526_ (.A0(_05399_),
    .A1(\tag_array.tag0[10][17] ),
    .S(_05567_),
    .X(_01279_));
 sky130_fd_sc_hd__mux2_1 _09527_ (.A0(_05401_),
    .A1(\tag_array.tag0[10][18] ),
    .S(_05567_),
    .X(_01280_));
 sky130_fd_sc_hd__mux2_1 _09528_ (.A0(_05403_),
    .A1(\tag_array.tag0[10][19] ),
    .S(_05567_),
    .X(_01281_));
 sky130_fd_sc_hd__mux2_1 _09529_ (.A0(_05405_),
    .A1(\tag_array.tag0[10][20] ),
    .S(_05567_),
    .X(_01282_));
 sky130_fd_sc_hd__mux2_1 _09530_ (.A0(_05407_),
    .A1(\tag_array.tag0[10][21] ),
    .S(_05567_),
    .X(_01283_));
 sky130_fd_sc_hd__mux2_1 _09531_ (.A0(_05409_),
    .A1(\tag_array.tag0[10][22] ),
    .S(_05567_),
    .X(_01284_));
 sky130_fd_sc_hd__mux2_1 _09532_ (.A0(_05411_),
    .A1(\tag_array.tag0[10][23] ),
    .S(_05567_),
    .X(_01285_));
 sky130_fd_sc_hd__mux2_1 _09533_ (.A0(_05413_),
    .A1(\tag_array.tag0[10][24] ),
    .S(_05567_),
    .X(_01286_));
 sky130_fd_sc_hd__mux2_1 _09534_ (.A0(_05365_),
    .A1(\tag_array.tag0[0][0] ),
    .S(_05569_),
    .X(_01287_));
 sky130_fd_sc_hd__mux2_1 _09535_ (.A0(_05367_),
    .A1(\tag_array.tag0[0][1] ),
    .S(_05569_),
    .X(_01288_));
 sky130_fd_sc_hd__mux2_1 _09536_ (.A0(_05369_),
    .A1(\tag_array.tag0[0][2] ),
    .S(_05569_),
    .X(_01289_));
 sky130_fd_sc_hd__mux2_1 _09537_ (.A0(_05371_),
    .A1(\tag_array.tag0[0][3] ),
    .S(_05569_),
    .X(_01290_));
 sky130_fd_sc_hd__mux2_1 _09538_ (.A0(_05373_),
    .A1(\tag_array.tag0[0][4] ),
    .S(_05569_),
    .X(_01291_));
 sky130_fd_sc_hd__mux2_1 _09539_ (.A0(_05375_),
    .A1(\tag_array.tag0[0][5] ),
    .S(_05569_),
    .X(_01292_));
 sky130_fd_sc_hd__mux2_1 _09540_ (.A0(_05377_),
    .A1(\tag_array.tag0[0][6] ),
    .S(_05569_),
    .X(_01293_));
 sky130_fd_sc_hd__mux2_1 _09541_ (.A0(_05379_),
    .A1(\tag_array.tag0[0][7] ),
    .S(_05569_),
    .X(_01294_));
 sky130_fd_sc_hd__mux2_1 _09542_ (.A0(_05381_),
    .A1(\tag_array.tag0[0][8] ),
    .S(_05569_),
    .X(_01295_));
 sky130_fd_sc_hd__mux2_1 _09543_ (.A0(_05383_),
    .A1(\tag_array.tag0[0][9] ),
    .S(_05569_),
    .X(_01296_));
 sky130_fd_sc_hd__mux2_1 _09544_ (.A0(_05385_),
    .A1(\tag_array.tag0[0][10] ),
    .S(_05569_),
    .X(_01297_));
 sky130_fd_sc_hd__mux2_1 _09545_ (.A0(_05387_),
    .A1(\tag_array.tag0[0][11] ),
    .S(_05569_),
    .X(_01298_));
 sky130_fd_sc_hd__mux2_1 _09546_ (.A0(_05389_),
    .A1(\tag_array.tag0[0][12] ),
    .S(_05569_),
    .X(_01299_));
 sky130_fd_sc_hd__mux2_1 _09547_ (.A0(_05391_),
    .A1(\tag_array.tag0[0][13] ),
    .S(_05569_),
    .X(_01300_));
 sky130_fd_sc_hd__mux2_1 _09548_ (.A0(_05393_),
    .A1(\tag_array.tag0[0][14] ),
    .S(_05569_),
    .X(_01301_));
 sky130_fd_sc_hd__mux2_1 _09549_ (.A0(_05395_),
    .A1(\tag_array.tag0[0][15] ),
    .S(_05569_),
    .X(_01302_));
 sky130_fd_sc_hd__mux2_1 _09550_ (.A0(_05397_),
    .A1(\tag_array.tag0[0][16] ),
    .S(_05569_),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_1 _09551_ (.A0(_05399_),
    .A1(\tag_array.tag0[0][17] ),
    .S(_05569_),
    .X(_01304_));
 sky130_fd_sc_hd__mux2_1 _09552_ (.A0(_05401_),
    .A1(\tag_array.tag0[0][18] ),
    .S(_05569_),
    .X(_01305_));
 sky130_fd_sc_hd__mux2_1 _09553_ (.A0(_05403_),
    .A1(\tag_array.tag0[0][19] ),
    .S(_05569_),
    .X(_01306_));
 sky130_fd_sc_hd__mux2_1 _09554_ (.A0(_05405_),
    .A1(\tag_array.tag0[0][20] ),
    .S(_05569_),
    .X(_01307_));
 sky130_fd_sc_hd__mux2_1 _09555_ (.A0(_05407_),
    .A1(\tag_array.tag0[0][21] ),
    .S(_05569_),
    .X(_01308_));
 sky130_fd_sc_hd__mux2_1 _09556_ (.A0(_05409_),
    .A1(\tag_array.tag0[0][22] ),
    .S(_05569_),
    .X(_01309_));
 sky130_fd_sc_hd__mux2_1 _09557_ (.A0(_05411_),
    .A1(\tag_array.tag0[0][23] ),
    .S(_05569_),
    .X(_01310_));
 sky130_fd_sc_hd__mux2_1 _09558_ (.A0(_05413_),
    .A1(\tag_array.tag0[0][24] ),
    .S(_05569_),
    .X(_01311_));
 sky130_fd_sc_hd__or2_2 _09559_ (.A(_05414_),
    .B(_05595_),
    .X(_03124_));
 sky130_fd_sc_hd__mux2_1 _09560_ (.A0(_05420_),
    .A1(\data_array.data0[15][0] ),
    .S(_03124_),
    .X(_01312_));
 sky130_fd_sc_hd__mux2_1 _09561_ (.A0(_05422_),
    .A1(\data_array.data0[15][1] ),
    .S(_03124_),
    .X(_01313_));
 sky130_fd_sc_hd__mux2_1 _09562_ (.A0(_05424_),
    .A1(\data_array.data0[15][2] ),
    .S(_03124_),
    .X(_01314_));
 sky130_fd_sc_hd__mux2_1 _09563_ (.A0(_05426_),
    .A1(\data_array.data0[15][3] ),
    .S(_03124_),
    .X(_01315_));
 sky130_fd_sc_hd__mux2_1 _09564_ (.A0(_05428_),
    .A1(\data_array.data0[15][4] ),
    .S(_03124_),
    .X(_01316_));
 sky130_fd_sc_hd__mux2_1 _09565_ (.A0(_05430_),
    .A1(\data_array.data0[15][5] ),
    .S(_03124_),
    .X(_01317_));
 sky130_fd_sc_hd__mux2_1 _09566_ (.A0(_05432_),
    .A1(\data_array.data0[15][6] ),
    .S(_03124_),
    .X(_01318_));
 sky130_fd_sc_hd__mux2_1 _09567_ (.A0(_05434_),
    .A1(\data_array.data0[15][7] ),
    .S(_03124_),
    .X(_01319_));
 sky130_fd_sc_hd__mux2_1 _09568_ (.A0(_05436_),
    .A1(\data_array.data0[15][8] ),
    .S(_03124_),
    .X(_01320_));
 sky130_fd_sc_hd__mux2_1 _09569_ (.A0(_05438_),
    .A1(\data_array.data0[15][9] ),
    .S(_03124_),
    .X(_01321_));
 sky130_fd_sc_hd__mux2_1 _09570_ (.A0(_05440_),
    .A1(\data_array.data0[15][10] ),
    .S(_03124_),
    .X(_01322_));
 sky130_fd_sc_hd__mux2_1 _09571_ (.A0(_05442_),
    .A1(\data_array.data0[15][11] ),
    .S(_03124_),
    .X(_01323_));
 sky130_fd_sc_hd__mux2_1 _09572_ (.A0(_05444_),
    .A1(\data_array.data0[15][12] ),
    .S(_03124_),
    .X(_01324_));
 sky130_fd_sc_hd__mux2_1 _09573_ (.A0(_05446_),
    .A1(\data_array.data0[15][13] ),
    .S(_03124_),
    .X(_01325_));
 sky130_fd_sc_hd__mux2_1 _09574_ (.A0(_05448_),
    .A1(\data_array.data0[15][14] ),
    .S(_03124_),
    .X(_01326_));
 sky130_fd_sc_hd__mux2_1 _09575_ (.A0(_05450_),
    .A1(\data_array.data0[15][15] ),
    .S(_03124_),
    .X(_01327_));
 sky130_fd_sc_hd__mux2_1 _09576_ (.A0(_05452_),
    .A1(\data_array.data0[15][16] ),
    .S(_03124_),
    .X(_01328_));
 sky130_fd_sc_hd__mux2_1 _09577_ (.A0(_05454_),
    .A1(\data_array.data0[15][17] ),
    .S(_03124_),
    .X(_01329_));
 sky130_fd_sc_hd__mux2_1 _09578_ (.A0(_05456_),
    .A1(\data_array.data0[15][18] ),
    .S(_03124_),
    .X(_01330_));
 sky130_fd_sc_hd__mux2_1 _09579_ (.A0(_05458_),
    .A1(\data_array.data0[15][19] ),
    .S(_03124_),
    .X(_01331_));
 sky130_fd_sc_hd__mux2_1 _09580_ (.A0(_05460_),
    .A1(\data_array.data0[15][20] ),
    .S(_03124_),
    .X(_01332_));
 sky130_fd_sc_hd__mux2_1 _09581_ (.A0(_05462_),
    .A1(\data_array.data0[15][21] ),
    .S(_03124_),
    .X(_01333_));
 sky130_fd_sc_hd__mux2_1 _09582_ (.A0(_05464_),
    .A1(\data_array.data0[15][22] ),
    .S(_03124_),
    .X(_01334_));
 sky130_fd_sc_hd__mux2_1 _09583_ (.A0(_05466_),
    .A1(\data_array.data0[15][23] ),
    .S(_03124_),
    .X(_01335_));
 sky130_fd_sc_hd__mux2_1 _09584_ (.A0(_05468_),
    .A1(\data_array.data0[15][24] ),
    .S(_03124_),
    .X(_01336_));
 sky130_fd_sc_hd__mux2_1 _09585_ (.A0(_05470_),
    .A1(\data_array.data0[15][25] ),
    .S(_03124_),
    .X(_01337_));
 sky130_fd_sc_hd__mux2_1 _09586_ (.A0(_05472_),
    .A1(\data_array.data0[15][26] ),
    .S(_03124_),
    .X(_01338_));
 sky130_fd_sc_hd__mux2_1 _09587_ (.A0(_05474_),
    .A1(\data_array.data0[15][27] ),
    .S(_03124_),
    .X(_01339_));
 sky130_fd_sc_hd__mux2_1 _09588_ (.A0(_05476_),
    .A1(\data_array.data0[15][28] ),
    .S(_03124_),
    .X(_01340_));
 sky130_fd_sc_hd__mux2_1 _09589_ (.A0(_05478_),
    .A1(\data_array.data0[15][29] ),
    .S(_03124_),
    .X(_01341_));
 sky130_fd_sc_hd__mux2_1 _09590_ (.A0(_05480_),
    .A1(\data_array.data0[15][30] ),
    .S(_03124_),
    .X(_01342_));
 sky130_fd_sc_hd__mux2_1 _09591_ (.A0(_05482_),
    .A1(\data_array.data0[15][31] ),
    .S(_03124_),
    .X(_01343_));
 sky130_fd_sc_hd__mux2_1 _09592_ (.A0(_05484_),
    .A1(\data_array.data0[15][32] ),
    .S(_03124_),
    .X(_01344_));
 sky130_fd_sc_hd__mux2_1 _09593_ (.A0(_05486_),
    .A1(\data_array.data0[15][33] ),
    .S(_03124_),
    .X(_01345_));
 sky130_fd_sc_hd__mux2_1 _09594_ (.A0(_05488_),
    .A1(\data_array.data0[15][34] ),
    .S(_03124_),
    .X(_01346_));
 sky130_fd_sc_hd__mux2_1 _09595_ (.A0(_05490_),
    .A1(\data_array.data0[15][35] ),
    .S(_03124_),
    .X(_01347_));
 sky130_fd_sc_hd__mux2_1 _09596_ (.A0(_05492_),
    .A1(\data_array.data0[15][36] ),
    .S(_03124_),
    .X(_01348_));
 sky130_fd_sc_hd__mux2_1 _09597_ (.A0(_05494_),
    .A1(\data_array.data0[15][37] ),
    .S(_03124_),
    .X(_01349_));
 sky130_fd_sc_hd__mux2_1 _09598_ (.A0(_05496_),
    .A1(\data_array.data0[15][38] ),
    .S(_03124_),
    .X(_01350_));
 sky130_fd_sc_hd__mux2_1 _09599_ (.A0(_05498_),
    .A1(\data_array.data0[15][39] ),
    .S(_03124_),
    .X(_01351_));
 sky130_fd_sc_hd__mux2_1 _09600_ (.A0(_05500_),
    .A1(\data_array.data0[15][40] ),
    .S(_03124_),
    .X(_01352_));
 sky130_fd_sc_hd__mux2_1 _09601_ (.A0(_05502_),
    .A1(\data_array.data0[15][41] ),
    .S(_03124_),
    .X(_01353_));
 sky130_fd_sc_hd__mux2_1 _09602_ (.A0(_05504_),
    .A1(\data_array.data0[15][42] ),
    .S(_03124_),
    .X(_01354_));
 sky130_fd_sc_hd__mux2_1 _09603_ (.A0(_05506_),
    .A1(\data_array.data0[15][43] ),
    .S(_03124_),
    .X(_01355_));
 sky130_fd_sc_hd__mux2_1 _09604_ (.A0(_05508_),
    .A1(\data_array.data0[15][44] ),
    .S(_03124_),
    .X(_01356_));
 sky130_fd_sc_hd__mux2_1 _09605_ (.A0(_05510_),
    .A1(\data_array.data0[15][45] ),
    .S(_03124_),
    .X(_01357_));
 sky130_fd_sc_hd__mux2_1 _09606_ (.A0(_05512_),
    .A1(\data_array.data0[15][46] ),
    .S(_03124_),
    .X(_01358_));
 sky130_fd_sc_hd__mux2_1 _09607_ (.A0(_05514_),
    .A1(\data_array.data0[15][47] ),
    .S(_03124_),
    .X(_01359_));
 sky130_fd_sc_hd__mux2_1 _09608_ (.A0(_05516_),
    .A1(\data_array.data0[15][48] ),
    .S(_03124_),
    .X(_01360_));
 sky130_fd_sc_hd__mux2_1 _09609_ (.A0(_05518_),
    .A1(\data_array.data0[15][49] ),
    .S(_03124_),
    .X(_01361_));
 sky130_fd_sc_hd__mux2_1 _09610_ (.A0(_05520_),
    .A1(\data_array.data0[15][50] ),
    .S(_03124_),
    .X(_01362_));
 sky130_fd_sc_hd__mux2_1 _09611_ (.A0(_05522_),
    .A1(\data_array.data0[15][51] ),
    .S(_03124_),
    .X(_01363_));
 sky130_fd_sc_hd__mux2_1 _09612_ (.A0(_05524_),
    .A1(\data_array.data0[15][52] ),
    .S(_03124_),
    .X(_01364_));
 sky130_fd_sc_hd__mux2_1 _09613_ (.A0(_05526_),
    .A1(\data_array.data0[15][53] ),
    .S(_03124_),
    .X(_01365_));
 sky130_fd_sc_hd__mux2_1 _09614_ (.A0(_05528_),
    .A1(\data_array.data0[15][54] ),
    .S(_03124_),
    .X(_01366_));
 sky130_fd_sc_hd__mux2_1 _09615_ (.A0(_05530_),
    .A1(\data_array.data0[15][55] ),
    .S(_03124_),
    .X(_01367_));
 sky130_fd_sc_hd__mux2_1 _09616_ (.A0(_05532_),
    .A1(\data_array.data0[15][56] ),
    .S(_03124_),
    .X(_01368_));
 sky130_fd_sc_hd__mux2_1 _09617_ (.A0(_05534_),
    .A1(\data_array.data0[15][57] ),
    .S(_03124_),
    .X(_01369_));
 sky130_fd_sc_hd__mux2_1 _09618_ (.A0(_05536_),
    .A1(\data_array.data0[15][58] ),
    .S(_03124_),
    .X(_01370_));
 sky130_fd_sc_hd__mux2_1 _09619_ (.A0(_05538_),
    .A1(\data_array.data0[15][59] ),
    .S(_03124_),
    .X(_01371_));
 sky130_fd_sc_hd__mux2_1 _09620_ (.A0(_05540_),
    .A1(\data_array.data0[15][60] ),
    .S(_03124_),
    .X(_01372_));
 sky130_fd_sc_hd__mux2_1 _09621_ (.A0(_05542_),
    .A1(\data_array.data0[15][61] ),
    .S(_03124_),
    .X(_01373_));
 sky130_fd_sc_hd__mux2_1 _09622_ (.A0(_05544_),
    .A1(\data_array.data0[15][62] ),
    .S(_03124_),
    .X(_01374_));
 sky130_fd_sc_hd__mux2_1 _09623_ (.A0(_05546_),
    .A1(\data_array.data0[15][63] ),
    .S(_03124_),
    .X(_01375_));
 sky130_fd_sc_hd__mux2_1 _09624_ (.A0(_05365_),
    .A1(\tag_array.tag0[8][0] ),
    .S(_05571_),
    .X(_01376_));
 sky130_fd_sc_hd__mux2_1 _09625_ (.A0(_05367_),
    .A1(\tag_array.tag0[8][1] ),
    .S(_05571_),
    .X(_01377_));
 sky130_fd_sc_hd__mux2_1 _09626_ (.A0(_05369_),
    .A1(\tag_array.tag0[8][2] ),
    .S(_05571_),
    .X(_01378_));
 sky130_fd_sc_hd__mux2_1 _09627_ (.A0(_05371_),
    .A1(\tag_array.tag0[8][3] ),
    .S(_05571_),
    .X(_01379_));
 sky130_fd_sc_hd__mux2_1 _09628_ (.A0(_05373_),
    .A1(\tag_array.tag0[8][4] ),
    .S(_05571_),
    .X(_01380_));
 sky130_fd_sc_hd__mux2_1 _09629_ (.A0(_05375_),
    .A1(\tag_array.tag0[8][5] ),
    .S(_05571_),
    .X(_01381_));
 sky130_fd_sc_hd__mux2_1 _09630_ (.A0(_05377_),
    .A1(\tag_array.tag0[8][6] ),
    .S(_05571_),
    .X(_01382_));
 sky130_fd_sc_hd__mux2_1 _09631_ (.A0(_05379_),
    .A1(\tag_array.tag0[8][7] ),
    .S(_05571_),
    .X(_01383_));
 sky130_fd_sc_hd__mux2_1 _09632_ (.A0(_05381_),
    .A1(\tag_array.tag0[8][8] ),
    .S(_05571_),
    .X(_01384_));
 sky130_fd_sc_hd__mux2_1 _09633_ (.A0(_05383_),
    .A1(\tag_array.tag0[8][9] ),
    .S(_05571_),
    .X(_01385_));
 sky130_fd_sc_hd__mux2_1 _09634_ (.A0(_05385_),
    .A1(\tag_array.tag0[8][10] ),
    .S(_05571_),
    .X(_01386_));
 sky130_fd_sc_hd__mux2_1 _09635_ (.A0(_05387_),
    .A1(\tag_array.tag0[8][11] ),
    .S(_05571_),
    .X(_01387_));
 sky130_fd_sc_hd__mux2_1 _09636_ (.A0(_05389_),
    .A1(\tag_array.tag0[8][12] ),
    .S(_05571_),
    .X(_01388_));
 sky130_fd_sc_hd__mux2_1 _09637_ (.A0(_05391_),
    .A1(\tag_array.tag0[8][13] ),
    .S(_05571_),
    .X(_01389_));
 sky130_fd_sc_hd__mux2_1 _09638_ (.A0(_05393_),
    .A1(\tag_array.tag0[8][14] ),
    .S(_05571_),
    .X(_01390_));
 sky130_fd_sc_hd__mux2_1 _09639_ (.A0(_05395_),
    .A1(\tag_array.tag0[8][15] ),
    .S(_05571_),
    .X(_01391_));
 sky130_fd_sc_hd__mux2_1 _09640_ (.A0(_05397_),
    .A1(\tag_array.tag0[8][16] ),
    .S(_05571_),
    .X(_01392_));
 sky130_fd_sc_hd__mux2_1 _09641_ (.A0(_05399_),
    .A1(\tag_array.tag0[8][17] ),
    .S(_05571_),
    .X(_01393_));
 sky130_fd_sc_hd__mux2_1 _09642_ (.A0(_05401_),
    .A1(\tag_array.tag0[8][18] ),
    .S(_05571_),
    .X(_01394_));
 sky130_fd_sc_hd__mux2_1 _09643_ (.A0(_05403_),
    .A1(\tag_array.tag0[8][19] ),
    .S(_05571_),
    .X(_01395_));
 sky130_fd_sc_hd__mux2_1 _09644_ (.A0(_05405_),
    .A1(\tag_array.tag0[8][20] ),
    .S(_05571_),
    .X(_01396_));
 sky130_fd_sc_hd__mux2_1 _09645_ (.A0(_05407_),
    .A1(\tag_array.tag0[8][21] ),
    .S(_05571_),
    .X(_01397_));
 sky130_fd_sc_hd__mux2_1 _09646_ (.A0(_05409_),
    .A1(\tag_array.tag0[8][22] ),
    .S(_05571_),
    .X(_01398_));
 sky130_fd_sc_hd__mux2_1 _09647_ (.A0(_05411_),
    .A1(\tag_array.tag0[8][23] ),
    .S(_05571_),
    .X(_01399_));
 sky130_fd_sc_hd__mux2_1 _09648_ (.A0(_05413_),
    .A1(\tag_array.tag0[8][24] ),
    .S(_05571_),
    .X(_01400_));
 sky130_fd_sc_hd__mux2_1 _09649_ (.A0(_05365_),
    .A1(\tag_array.tag0[7][0] ),
    .S(_05573_),
    .X(_01401_));
 sky130_fd_sc_hd__mux2_1 _09650_ (.A0(_05367_),
    .A1(\tag_array.tag0[7][1] ),
    .S(_05573_),
    .X(_01402_));
 sky130_fd_sc_hd__mux2_1 _09651_ (.A0(_05369_),
    .A1(\tag_array.tag0[7][2] ),
    .S(_05573_),
    .X(_01403_));
 sky130_fd_sc_hd__mux2_1 _09652_ (.A0(_05371_),
    .A1(\tag_array.tag0[7][3] ),
    .S(_05573_),
    .X(_01404_));
 sky130_fd_sc_hd__mux2_1 _09653_ (.A0(_05373_),
    .A1(\tag_array.tag0[7][4] ),
    .S(_05573_),
    .X(_01405_));
 sky130_fd_sc_hd__mux2_1 _09654_ (.A0(_05375_),
    .A1(\tag_array.tag0[7][5] ),
    .S(_05573_),
    .X(_01406_));
 sky130_fd_sc_hd__mux2_1 _09655_ (.A0(_05377_),
    .A1(\tag_array.tag0[7][6] ),
    .S(_05573_),
    .X(_01407_));
 sky130_fd_sc_hd__mux2_1 _09656_ (.A0(_05379_),
    .A1(\tag_array.tag0[7][7] ),
    .S(_05573_),
    .X(_01408_));
 sky130_fd_sc_hd__mux2_1 _09657_ (.A0(_05381_),
    .A1(\tag_array.tag0[7][8] ),
    .S(_05573_),
    .X(_01409_));
 sky130_fd_sc_hd__mux2_1 _09658_ (.A0(_05383_),
    .A1(\tag_array.tag0[7][9] ),
    .S(_05573_),
    .X(_01410_));
 sky130_fd_sc_hd__mux2_1 _09659_ (.A0(_05385_),
    .A1(\tag_array.tag0[7][10] ),
    .S(_05573_),
    .X(_01411_));
 sky130_fd_sc_hd__mux2_1 _09660_ (.A0(_05387_),
    .A1(\tag_array.tag0[7][11] ),
    .S(_05573_),
    .X(_01412_));
 sky130_fd_sc_hd__mux2_1 _09661_ (.A0(_05389_),
    .A1(\tag_array.tag0[7][12] ),
    .S(_05573_),
    .X(_01413_));
 sky130_fd_sc_hd__mux2_1 _09662_ (.A0(_05391_),
    .A1(\tag_array.tag0[7][13] ),
    .S(_05573_),
    .X(_01414_));
 sky130_fd_sc_hd__mux2_1 _09663_ (.A0(_05393_),
    .A1(\tag_array.tag0[7][14] ),
    .S(_05573_),
    .X(_01415_));
 sky130_fd_sc_hd__mux2_1 _09664_ (.A0(_05395_),
    .A1(\tag_array.tag0[7][15] ),
    .S(_05573_),
    .X(_01416_));
 sky130_fd_sc_hd__mux2_1 _09665_ (.A0(_05397_),
    .A1(\tag_array.tag0[7][16] ),
    .S(_05573_),
    .X(_01417_));
 sky130_fd_sc_hd__mux2_1 _09666_ (.A0(_05399_),
    .A1(\tag_array.tag0[7][17] ),
    .S(_05573_),
    .X(_01418_));
 sky130_fd_sc_hd__mux2_1 _09667_ (.A0(_05401_),
    .A1(\tag_array.tag0[7][18] ),
    .S(_05573_),
    .X(_01419_));
 sky130_fd_sc_hd__mux2_1 _09668_ (.A0(_05403_),
    .A1(\tag_array.tag0[7][19] ),
    .S(_05573_),
    .X(_01420_));
 sky130_fd_sc_hd__mux2_1 _09669_ (.A0(_05405_),
    .A1(\tag_array.tag0[7][20] ),
    .S(_05573_),
    .X(_01421_));
 sky130_fd_sc_hd__mux2_1 _09670_ (.A0(_05407_),
    .A1(\tag_array.tag0[7][21] ),
    .S(_05573_),
    .X(_01422_));
 sky130_fd_sc_hd__mux2_1 _09671_ (.A0(_05409_),
    .A1(\tag_array.tag0[7][22] ),
    .S(_05573_),
    .X(_01423_));
 sky130_fd_sc_hd__mux2_1 _09672_ (.A0(_05411_),
    .A1(\tag_array.tag0[7][23] ),
    .S(_05573_),
    .X(_01424_));
 sky130_fd_sc_hd__mux2_1 _09673_ (.A0(_05413_),
    .A1(\tag_array.tag0[7][24] ),
    .S(_05573_),
    .X(_01425_));
 sky130_fd_sc_hd__mux2_1 _09674_ (.A0(_05365_),
    .A1(\tag_array.tag0[5][0] ),
    .S(_05579_),
    .X(_01426_));
 sky130_fd_sc_hd__mux2_1 _09675_ (.A0(_05367_),
    .A1(\tag_array.tag0[5][1] ),
    .S(_05579_),
    .X(_01427_));
 sky130_fd_sc_hd__mux2_1 _09676_ (.A0(_05369_),
    .A1(\tag_array.tag0[5][2] ),
    .S(_05579_),
    .X(_01428_));
 sky130_fd_sc_hd__mux2_1 _09677_ (.A0(_05371_),
    .A1(\tag_array.tag0[5][3] ),
    .S(_05579_),
    .X(_01429_));
 sky130_fd_sc_hd__mux2_1 _09678_ (.A0(_05373_),
    .A1(\tag_array.tag0[5][4] ),
    .S(_05579_),
    .X(_01430_));
 sky130_fd_sc_hd__mux2_1 _09679_ (.A0(_05375_),
    .A1(\tag_array.tag0[5][5] ),
    .S(_05579_),
    .X(_01431_));
 sky130_fd_sc_hd__mux2_1 _09680_ (.A0(_05377_),
    .A1(\tag_array.tag0[5][6] ),
    .S(_05579_),
    .X(_01432_));
 sky130_fd_sc_hd__mux2_1 _09681_ (.A0(_05379_),
    .A1(\tag_array.tag0[5][7] ),
    .S(_05579_),
    .X(_01433_));
 sky130_fd_sc_hd__mux2_1 _09682_ (.A0(_05381_),
    .A1(\tag_array.tag0[5][8] ),
    .S(_05579_),
    .X(_01434_));
 sky130_fd_sc_hd__mux2_1 _09683_ (.A0(_05383_),
    .A1(\tag_array.tag0[5][9] ),
    .S(_05579_),
    .X(_01435_));
 sky130_fd_sc_hd__mux2_1 _09684_ (.A0(_05385_),
    .A1(\tag_array.tag0[5][10] ),
    .S(_05579_),
    .X(_01436_));
 sky130_fd_sc_hd__mux2_1 _09685_ (.A0(_05387_),
    .A1(\tag_array.tag0[5][11] ),
    .S(_05579_),
    .X(_01437_));
 sky130_fd_sc_hd__mux2_1 _09686_ (.A0(_05389_),
    .A1(\tag_array.tag0[5][12] ),
    .S(_05579_),
    .X(_01438_));
 sky130_fd_sc_hd__mux2_1 _09687_ (.A0(_05391_),
    .A1(\tag_array.tag0[5][13] ),
    .S(_05579_),
    .X(_01439_));
 sky130_fd_sc_hd__mux2_1 _09688_ (.A0(_05393_),
    .A1(\tag_array.tag0[5][14] ),
    .S(_05579_),
    .X(_01440_));
 sky130_fd_sc_hd__mux2_1 _09689_ (.A0(_05395_),
    .A1(\tag_array.tag0[5][15] ),
    .S(_05579_),
    .X(_01441_));
 sky130_fd_sc_hd__mux2_1 _09690_ (.A0(_05397_),
    .A1(\tag_array.tag0[5][16] ),
    .S(_05579_),
    .X(_01442_));
 sky130_fd_sc_hd__mux2_1 _09691_ (.A0(_05399_),
    .A1(\tag_array.tag0[5][17] ),
    .S(_05579_),
    .X(_01443_));
 sky130_fd_sc_hd__mux2_1 _09692_ (.A0(_05401_),
    .A1(\tag_array.tag0[5][18] ),
    .S(_05579_),
    .X(_01444_));
 sky130_fd_sc_hd__mux2_1 _09693_ (.A0(_05403_),
    .A1(\tag_array.tag0[5][19] ),
    .S(_05579_),
    .X(_01445_));
 sky130_fd_sc_hd__mux2_1 _09694_ (.A0(_05405_),
    .A1(\tag_array.tag0[5][20] ),
    .S(_05579_),
    .X(_01446_));
 sky130_fd_sc_hd__mux2_1 _09695_ (.A0(_05407_),
    .A1(\tag_array.tag0[5][21] ),
    .S(_05579_),
    .X(_01447_));
 sky130_fd_sc_hd__mux2_1 _09696_ (.A0(_05409_),
    .A1(\tag_array.tag0[5][22] ),
    .S(_05579_),
    .X(_01448_));
 sky130_fd_sc_hd__mux2_1 _09697_ (.A0(_05411_),
    .A1(\tag_array.tag0[5][23] ),
    .S(_05579_),
    .X(_01449_));
 sky130_fd_sc_hd__mux2_1 _09698_ (.A0(_05413_),
    .A1(\tag_array.tag0[5][24] ),
    .S(_05579_),
    .X(_01450_));
 sky130_fd_sc_hd__mux2_1 _09699_ (.A0(_05365_),
    .A1(\tag_array.tag0[6][0] ),
    .S(_05576_),
    .X(_01451_));
 sky130_fd_sc_hd__mux2_1 _09700_ (.A0(_05367_),
    .A1(\tag_array.tag0[6][1] ),
    .S(_05576_),
    .X(_01452_));
 sky130_fd_sc_hd__mux2_1 _09701_ (.A0(_05369_),
    .A1(\tag_array.tag0[6][2] ),
    .S(_05576_),
    .X(_01453_));
 sky130_fd_sc_hd__mux2_1 _09702_ (.A0(_05371_),
    .A1(\tag_array.tag0[6][3] ),
    .S(_05576_),
    .X(_01454_));
 sky130_fd_sc_hd__mux2_1 _09703_ (.A0(_05373_),
    .A1(\tag_array.tag0[6][4] ),
    .S(_05576_),
    .X(_01455_));
 sky130_fd_sc_hd__mux2_1 _09704_ (.A0(_05375_),
    .A1(\tag_array.tag0[6][5] ),
    .S(_05576_),
    .X(_01456_));
 sky130_fd_sc_hd__mux2_1 _09705_ (.A0(_05377_),
    .A1(\tag_array.tag0[6][6] ),
    .S(_05576_),
    .X(_01457_));
 sky130_fd_sc_hd__mux2_1 _09706_ (.A0(_05379_),
    .A1(\tag_array.tag0[6][7] ),
    .S(_05576_),
    .X(_01458_));
 sky130_fd_sc_hd__mux2_1 _09707_ (.A0(_05381_),
    .A1(\tag_array.tag0[6][8] ),
    .S(_05576_),
    .X(_01459_));
 sky130_fd_sc_hd__mux2_1 _09708_ (.A0(_05383_),
    .A1(\tag_array.tag0[6][9] ),
    .S(_05576_),
    .X(_01460_));
 sky130_fd_sc_hd__mux2_1 _09709_ (.A0(_05385_),
    .A1(\tag_array.tag0[6][10] ),
    .S(_05576_),
    .X(_01461_));
 sky130_fd_sc_hd__mux2_1 _09710_ (.A0(_05387_),
    .A1(\tag_array.tag0[6][11] ),
    .S(_05576_),
    .X(_01462_));
 sky130_fd_sc_hd__mux2_1 _09711_ (.A0(_05389_),
    .A1(\tag_array.tag0[6][12] ),
    .S(_05576_),
    .X(_01463_));
 sky130_fd_sc_hd__mux2_1 _09712_ (.A0(_05391_),
    .A1(\tag_array.tag0[6][13] ),
    .S(_05576_),
    .X(_01464_));
 sky130_fd_sc_hd__mux2_1 _09713_ (.A0(_05393_),
    .A1(\tag_array.tag0[6][14] ),
    .S(_05576_),
    .X(_01465_));
 sky130_fd_sc_hd__mux2_1 _09714_ (.A0(_05395_),
    .A1(\tag_array.tag0[6][15] ),
    .S(_05576_),
    .X(_01466_));
 sky130_fd_sc_hd__mux2_1 _09715_ (.A0(_05397_),
    .A1(\tag_array.tag0[6][16] ),
    .S(_05576_),
    .X(_01467_));
 sky130_fd_sc_hd__mux2_1 _09716_ (.A0(_05399_),
    .A1(\tag_array.tag0[6][17] ),
    .S(_05576_),
    .X(_01468_));
 sky130_fd_sc_hd__mux2_1 _09717_ (.A0(_05401_),
    .A1(\tag_array.tag0[6][18] ),
    .S(_05576_),
    .X(_01469_));
 sky130_fd_sc_hd__mux2_1 _09718_ (.A0(_05403_),
    .A1(\tag_array.tag0[6][19] ),
    .S(_05576_),
    .X(_01470_));
 sky130_fd_sc_hd__mux2_1 _09719_ (.A0(_05405_),
    .A1(\tag_array.tag0[6][20] ),
    .S(_05576_),
    .X(_01471_));
 sky130_fd_sc_hd__mux2_1 _09720_ (.A0(_05407_),
    .A1(\tag_array.tag0[6][21] ),
    .S(_05576_),
    .X(_01472_));
 sky130_fd_sc_hd__mux2_1 _09721_ (.A0(_05409_),
    .A1(\tag_array.tag0[6][22] ),
    .S(_05576_),
    .X(_01473_));
 sky130_fd_sc_hd__mux2_1 _09722_ (.A0(_05411_),
    .A1(\tag_array.tag0[6][23] ),
    .S(_05576_),
    .X(_01474_));
 sky130_fd_sc_hd__mux2_1 _09723_ (.A0(_05413_),
    .A1(\tag_array.tag0[6][24] ),
    .S(_05576_),
    .X(_01475_));
 sky130_fd_sc_hd__mux2_1 _09724_ (.A0(_05365_),
    .A1(\tag_array.tag1[10][0] ),
    .S(_05548_),
    .X(_01476_));
 sky130_fd_sc_hd__mux2_1 _09725_ (.A0(_05367_),
    .A1(\tag_array.tag1[10][1] ),
    .S(_05548_),
    .X(_01477_));
 sky130_fd_sc_hd__mux2_1 _09726_ (.A0(_05369_),
    .A1(\tag_array.tag1[10][2] ),
    .S(_05548_),
    .X(_01478_));
 sky130_fd_sc_hd__mux2_1 _09727_ (.A0(_05371_),
    .A1(\tag_array.tag1[10][3] ),
    .S(_05548_),
    .X(_01479_));
 sky130_fd_sc_hd__mux2_1 _09728_ (.A0(_05373_),
    .A1(\tag_array.tag1[10][4] ),
    .S(_05548_),
    .X(_01480_));
 sky130_fd_sc_hd__mux2_1 _09729_ (.A0(_05375_),
    .A1(\tag_array.tag1[10][5] ),
    .S(_05548_),
    .X(_01481_));
 sky130_fd_sc_hd__mux2_1 _09730_ (.A0(_05377_),
    .A1(\tag_array.tag1[10][6] ),
    .S(_05548_),
    .X(_01482_));
 sky130_fd_sc_hd__mux2_1 _09731_ (.A0(_05379_),
    .A1(\tag_array.tag1[10][7] ),
    .S(_05548_),
    .X(_01483_));
 sky130_fd_sc_hd__mux2_1 _09732_ (.A0(_05381_),
    .A1(\tag_array.tag1[10][8] ),
    .S(_05548_),
    .X(_01484_));
 sky130_fd_sc_hd__mux2_1 _09733_ (.A0(_05383_),
    .A1(\tag_array.tag1[10][9] ),
    .S(_05548_),
    .X(_01485_));
 sky130_fd_sc_hd__mux2_1 _09734_ (.A0(_05385_),
    .A1(\tag_array.tag1[10][10] ),
    .S(_05548_),
    .X(_01486_));
 sky130_fd_sc_hd__mux2_1 _09735_ (.A0(_05387_),
    .A1(\tag_array.tag1[10][11] ),
    .S(_05548_),
    .X(_01487_));
 sky130_fd_sc_hd__mux2_1 _09736_ (.A0(_05389_),
    .A1(\tag_array.tag1[10][12] ),
    .S(_05548_),
    .X(_01488_));
 sky130_fd_sc_hd__mux2_1 _09737_ (.A0(_05391_),
    .A1(\tag_array.tag1[10][13] ),
    .S(_05548_),
    .X(_01489_));
 sky130_fd_sc_hd__mux2_1 _09738_ (.A0(_05393_),
    .A1(\tag_array.tag1[10][14] ),
    .S(_05548_),
    .X(_01490_));
 sky130_fd_sc_hd__mux2_1 _09739_ (.A0(_05395_),
    .A1(\tag_array.tag1[10][15] ),
    .S(_05548_),
    .X(_01491_));
 sky130_fd_sc_hd__mux2_1 _09740_ (.A0(_05397_),
    .A1(\tag_array.tag1[10][16] ),
    .S(_05548_),
    .X(_01492_));
 sky130_fd_sc_hd__mux2_1 _09741_ (.A0(_05399_),
    .A1(\tag_array.tag1[10][17] ),
    .S(_05548_),
    .X(_01493_));
 sky130_fd_sc_hd__mux2_1 _09742_ (.A0(_05401_),
    .A1(\tag_array.tag1[10][18] ),
    .S(_05548_),
    .X(_01494_));
 sky130_fd_sc_hd__mux2_1 _09743_ (.A0(_05403_),
    .A1(\tag_array.tag1[10][19] ),
    .S(_05548_),
    .X(_01495_));
 sky130_fd_sc_hd__mux2_1 _09744_ (.A0(_05405_),
    .A1(\tag_array.tag1[10][20] ),
    .S(_05548_),
    .X(_01496_));
 sky130_fd_sc_hd__mux2_1 _09745_ (.A0(_05407_),
    .A1(\tag_array.tag1[10][21] ),
    .S(_05548_),
    .X(_01497_));
 sky130_fd_sc_hd__mux2_1 _09746_ (.A0(_05409_),
    .A1(\tag_array.tag1[10][22] ),
    .S(_05548_),
    .X(_01498_));
 sky130_fd_sc_hd__mux2_1 _09747_ (.A0(_05411_),
    .A1(\tag_array.tag1[10][23] ),
    .S(_05548_),
    .X(_01499_));
 sky130_fd_sc_hd__mux2_1 _09748_ (.A0(_05413_),
    .A1(\tag_array.tag1[10][24] ),
    .S(_05548_),
    .X(_01500_));
 sky130_fd_sc_hd__mux2_1 _09749_ (.A0(\tag_array.tag1[0][0] ),
    .A1(_05365_),
    .S(_05549_),
    .X(_01501_));
 sky130_fd_sc_hd__mux2_1 _09750_ (.A0(\tag_array.tag1[0][1] ),
    .A1(_05367_),
    .S(_05549_),
    .X(_01502_));
 sky130_fd_sc_hd__mux2_1 _09751_ (.A0(\tag_array.tag1[0][2] ),
    .A1(_05369_),
    .S(_05549_),
    .X(_01503_));
 sky130_fd_sc_hd__mux2_1 _09752_ (.A0(\tag_array.tag1[0][3] ),
    .A1(_05371_),
    .S(_05549_),
    .X(_01504_));
 sky130_fd_sc_hd__mux2_1 _09753_ (.A0(\tag_array.tag1[0][4] ),
    .A1(_05373_),
    .S(_05549_),
    .X(_01505_));
 sky130_fd_sc_hd__mux2_1 _09754_ (.A0(\tag_array.tag1[0][5] ),
    .A1(_05375_),
    .S(_05549_),
    .X(_01506_));
 sky130_fd_sc_hd__mux2_1 _09755_ (.A0(\tag_array.tag1[0][6] ),
    .A1(_05377_),
    .S(_05549_),
    .X(_01507_));
 sky130_fd_sc_hd__mux2_1 _09756_ (.A0(\tag_array.tag1[0][7] ),
    .A1(_05379_),
    .S(_05549_),
    .X(_01508_));
 sky130_fd_sc_hd__mux2_1 _09757_ (.A0(\tag_array.tag1[0][8] ),
    .A1(_05381_),
    .S(_05549_),
    .X(_01509_));
 sky130_fd_sc_hd__mux2_1 _09758_ (.A0(\tag_array.tag1[0][9] ),
    .A1(_05383_),
    .S(_05549_),
    .X(_01510_));
 sky130_fd_sc_hd__mux2_1 _09759_ (.A0(\tag_array.tag1[0][10] ),
    .A1(_05385_),
    .S(_05549_),
    .X(_01511_));
 sky130_fd_sc_hd__mux2_1 _09760_ (.A0(\tag_array.tag1[0][11] ),
    .A1(_05387_),
    .S(_05549_),
    .X(_01512_));
 sky130_fd_sc_hd__mux2_1 _09761_ (.A0(\tag_array.tag1[0][12] ),
    .A1(_05389_),
    .S(_05549_),
    .X(_01513_));
 sky130_fd_sc_hd__mux2_1 _09762_ (.A0(\tag_array.tag1[0][13] ),
    .A1(_05391_),
    .S(_05549_),
    .X(_01514_));
 sky130_fd_sc_hd__mux2_1 _09763_ (.A0(\tag_array.tag1[0][14] ),
    .A1(_05393_),
    .S(_05549_),
    .X(_01515_));
 sky130_fd_sc_hd__mux2_1 _09764_ (.A0(\tag_array.tag1[0][15] ),
    .A1(_05395_),
    .S(_05549_),
    .X(_01516_));
 sky130_fd_sc_hd__mux2_1 _09765_ (.A0(\tag_array.tag1[0][16] ),
    .A1(_05397_),
    .S(_05549_),
    .X(_01517_));
 sky130_fd_sc_hd__mux2_1 _09766_ (.A0(\tag_array.tag1[0][17] ),
    .A1(_05399_),
    .S(_05549_),
    .X(_01518_));
 sky130_fd_sc_hd__mux2_1 _09767_ (.A0(\tag_array.tag1[0][18] ),
    .A1(_05401_),
    .S(_05549_),
    .X(_01519_));
 sky130_fd_sc_hd__mux2_1 _09768_ (.A0(\tag_array.tag1[0][19] ),
    .A1(_05403_),
    .S(_05549_),
    .X(_01520_));
 sky130_fd_sc_hd__mux2_1 _09769_ (.A0(\tag_array.tag1[0][20] ),
    .A1(_05405_),
    .S(_05549_),
    .X(_01521_));
 sky130_fd_sc_hd__mux2_1 _09770_ (.A0(\tag_array.tag1[0][21] ),
    .A1(_05407_),
    .S(_05549_),
    .X(_01522_));
 sky130_fd_sc_hd__mux2_1 _09771_ (.A0(\tag_array.tag1[0][22] ),
    .A1(_05409_),
    .S(_05549_),
    .X(_01523_));
 sky130_fd_sc_hd__mux2_1 _09772_ (.A0(\tag_array.tag1[0][23] ),
    .A1(_05411_),
    .S(_05549_),
    .X(_01524_));
 sky130_fd_sc_hd__mux2_1 _09773_ (.A0(\tag_array.tag1[0][24] ),
    .A1(_05413_),
    .S(_05549_),
    .X(_01525_));
 sky130_fd_sc_hd__nand2_2 _09774_ (.A(_05415_),
    .B(_05561_),
    .Y(_03125_));
 sky130_fd_sc_hd__mux2_1 _09775_ (.A0(_05420_),
    .A1(\data_array.data0[12][0] ),
    .S(_03125_),
    .X(_01526_));
 sky130_fd_sc_hd__mux2_1 _09776_ (.A0(_05422_),
    .A1(\data_array.data0[12][1] ),
    .S(_03125_),
    .X(_01527_));
 sky130_fd_sc_hd__mux2_1 _09777_ (.A0(_05424_),
    .A1(\data_array.data0[12][2] ),
    .S(_03125_),
    .X(_01528_));
 sky130_fd_sc_hd__mux2_1 _09778_ (.A0(_05426_),
    .A1(\data_array.data0[12][3] ),
    .S(_03125_),
    .X(_01529_));
 sky130_fd_sc_hd__mux2_1 _09779_ (.A0(_05428_),
    .A1(\data_array.data0[12][4] ),
    .S(_03125_),
    .X(_01530_));
 sky130_fd_sc_hd__mux2_1 _09780_ (.A0(_05430_),
    .A1(\data_array.data0[12][5] ),
    .S(_03125_),
    .X(_01531_));
 sky130_fd_sc_hd__mux2_1 _09781_ (.A0(_05432_),
    .A1(\data_array.data0[12][6] ),
    .S(_03125_),
    .X(_01532_));
 sky130_fd_sc_hd__mux2_1 _09782_ (.A0(_05434_),
    .A1(\data_array.data0[12][7] ),
    .S(_03125_),
    .X(_01533_));
 sky130_fd_sc_hd__mux2_1 _09783_ (.A0(_05436_),
    .A1(\data_array.data0[12][8] ),
    .S(_03125_),
    .X(_01534_));
 sky130_fd_sc_hd__mux2_1 _09784_ (.A0(_05438_),
    .A1(\data_array.data0[12][9] ),
    .S(_03125_),
    .X(_01535_));
 sky130_fd_sc_hd__mux2_1 _09785_ (.A0(_05440_),
    .A1(\data_array.data0[12][10] ),
    .S(_03125_),
    .X(_01536_));
 sky130_fd_sc_hd__mux2_1 _09786_ (.A0(_05442_),
    .A1(\data_array.data0[12][11] ),
    .S(_03125_),
    .X(_01537_));
 sky130_fd_sc_hd__mux2_1 _09787_ (.A0(_05444_),
    .A1(\data_array.data0[12][12] ),
    .S(_03125_),
    .X(_01538_));
 sky130_fd_sc_hd__mux2_1 _09788_ (.A0(_05446_),
    .A1(\data_array.data0[12][13] ),
    .S(_03125_),
    .X(_01539_));
 sky130_fd_sc_hd__mux2_1 _09789_ (.A0(_05448_),
    .A1(\data_array.data0[12][14] ),
    .S(_03125_),
    .X(_01540_));
 sky130_fd_sc_hd__mux2_1 _09790_ (.A0(_05450_),
    .A1(\data_array.data0[12][15] ),
    .S(_03125_),
    .X(_01541_));
 sky130_fd_sc_hd__mux2_1 _09791_ (.A0(_05452_),
    .A1(\data_array.data0[12][16] ),
    .S(_03125_),
    .X(_01542_));
 sky130_fd_sc_hd__mux2_1 _09792_ (.A0(_05454_),
    .A1(\data_array.data0[12][17] ),
    .S(_03125_),
    .X(_01543_));
 sky130_fd_sc_hd__mux2_1 _09793_ (.A0(_05456_),
    .A1(\data_array.data0[12][18] ),
    .S(_03125_),
    .X(_01544_));
 sky130_fd_sc_hd__mux2_1 _09794_ (.A0(_05458_),
    .A1(\data_array.data0[12][19] ),
    .S(_03125_),
    .X(_01545_));
 sky130_fd_sc_hd__mux2_1 _09795_ (.A0(_05460_),
    .A1(\data_array.data0[12][20] ),
    .S(_03125_),
    .X(_01546_));
 sky130_fd_sc_hd__mux2_1 _09796_ (.A0(_05462_),
    .A1(\data_array.data0[12][21] ),
    .S(_03125_),
    .X(_01547_));
 sky130_fd_sc_hd__mux2_1 _09797_ (.A0(_05464_),
    .A1(\data_array.data0[12][22] ),
    .S(_03125_),
    .X(_01548_));
 sky130_fd_sc_hd__mux2_1 _09798_ (.A0(_05466_),
    .A1(\data_array.data0[12][23] ),
    .S(_03125_),
    .X(_01549_));
 sky130_fd_sc_hd__mux2_1 _09799_ (.A0(_05468_),
    .A1(\data_array.data0[12][24] ),
    .S(_03125_),
    .X(_01550_));
 sky130_fd_sc_hd__mux2_1 _09800_ (.A0(_05470_),
    .A1(\data_array.data0[12][25] ),
    .S(_03125_),
    .X(_01551_));
 sky130_fd_sc_hd__mux2_1 _09801_ (.A0(_05472_),
    .A1(\data_array.data0[12][26] ),
    .S(_03125_),
    .X(_01552_));
 sky130_fd_sc_hd__mux2_1 _09802_ (.A0(_05474_),
    .A1(\data_array.data0[12][27] ),
    .S(_03125_),
    .X(_01553_));
 sky130_fd_sc_hd__mux2_1 _09803_ (.A0(_05476_),
    .A1(\data_array.data0[12][28] ),
    .S(_03125_),
    .X(_01554_));
 sky130_fd_sc_hd__mux2_1 _09804_ (.A0(_05478_),
    .A1(\data_array.data0[12][29] ),
    .S(_03125_),
    .X(_01555_));
 sky130_fd_sc_hd__mux2_1 _09805_ (.A0(_05480_),
    .A1(\data_array.data0[12][30] ),
    .S(_03125_),
    .X(_01556_));
 sky130_fd_sc_hd__mux2_1 _09806_ (.A0(_05482_),
    .A1(\data_array.data0[12][31] ),
    .S(_03125_),
    .X(_01557_));
 sky130_fd_sc_hd__mux2_1 _09807_ (.A0(_05484_),
    .A1(\data_array.data0[12][32] ),
    .S(_03125_),
    .X(_01558_));
 sky130_fd_sc_hd__mux2_1 _09808_ (.A0(_05486_),
    .A1(\data_array.data0[12][33] ),
    .S(_03125_),
    .X(_01559_));
 sky130_fd_sc_hd__mux2_1 _09809_ (.A0(_05488_),
    .A1(\data_array.data0[12][34] ),
    .S(_03125_),
    .X(_01560_));
 sky130_fd_sc_hd__mux2_1 _09810_ (.A0(_05490_),
    .A1(\data_array.data0[12][35] ),
    .S(_03125_),
    .X(_01561_));
 sky130_fd_sc_hd__mux2_1 _09811_ (.A0(_05492_),
    .A1(\data_array.data0[12][36] ),
    .S(_03125_),
    .X(_01562_));
 sky130_fd_sc_hd__mux2_1 _09812_ (.A0(_05494_),
    .A1(\data_array.data0[12][37] ),
    .S(_03125_),
    .X(_01563_));
 sky130_fd_sc_hd__mux2_1 _09813_ (.A0(_05496_),
    .A1(\data_array.data0[12][38] ),
    .S(_03125_),
    .X(_01564_));
 sky130_fd_sc_hd__mux2_1 _09814_ (.A0(_05498_),
    .A1(\data_array.data0[12][39] ),
    .S(_03125_),
    .X(_01565_));
 sky130_fd_sc_hd__mux2_1 _09815_ (.A0(_05500_),
    .A1(\data_array.data0[12][40] ),
    .S(_03125_),
    .X(_01566_));
 sky130_fd_sc_hd__mux2_1 _09816_ (.A0(_05502_),
    .A1(\data_array.data0[12][41] ),
    .S(_03125_),
    .X(_01567_));
 sky130_fd_sc_hd__mux2_1 _09817_ (.A0(_05504_),
    .A1(\data_array.data0[12][42] ),
    .S(_03125_),
    .X(_01568_));
 sky130_fd_sc_hd__mux2_1 _09818_ (.A0(_05506_),
    .A1(\data_array.data0[12][43] ),
    .S(_03125_),
    .X(_01569_));
 sky130_fd_sc_hd__mux2_1 _09819_ (.A0(_05508_),
    .A1(\data_array.data0[12][44] ),
    .S(_03125_),
    .X(_01570_));
 sky130_fd_sc_hd__mux2_1 _09820_ (.A0(_05510_),
    .A1(\data_array.data0[12][45] ),
    .S(_03125_),
    .X(_01571_));
 sky130_fd_sc_hd__mux2_1 _09821_ (.A0(_05512_),
    .A1(\data_array.data0[12][46] ),
    .S(_03125_),
    .X(_01572_));
 sky130_fd_sc_hd__mux2_1 _09822_ (.A0(_05514_),
    .A1(\data_array.data0[12][47] ),
    .S(_03125_),
    .X(_01573_));
 sky130_fd_sc_hd__mux2_1 _09823_ (.A0(_05516_),
    .A1(\data_array.data0[12][48] ),
    .S(_03125_),
    .X(_01574_));
 sky130_fd_sc_hd__mux2_1 _09824_ (.A0(_05518_),
    .A1(\data_array.data0[12][49] ),
    .S(_03125_),
    .X(_01575_));
 sky130_fd_sc_hd__mux2_1 _09825_ (.A0(_05520_),
    .A1(\data_array.data0[12][50] ),
    .S(_03125_),
    .X(_01576_));
 sky130_fd_sc_hd__mux2_1 _09826_ (.A0(_05522_),
    .A1(\data_array.data0[12][51] ),
    .S(_03125_),
    .X(_01577_));
 sky130_fd_sc_hd__mux2_1 _09827_ (.A0(_05524_),
    .A1(\data_array.data0[12][52] ),
    .S(_03125_),
    .X(_01578_));
 sky130_fd_sc_hd__mux2_1 _09828_ (.A0(_05526_),
    .A1(\data_array.data0[12][53] ),
    .S(_03125_),
    .X(_01579_));
 sky130_fd_sc_hd__mux2_1 _09829_ (.A0(_05528_),
    .A1(\data_array.data0[12][54] ),
    .S(_03125_),
    .X(_01580_));
 sky130_fd_sc_hd__mux2_1 _09830_ (.A0(_05530_),
    .A1(\data_array.data0[12][55] ),
    .S(_03125_),
    .X(_01581_));
 sky130_fd_sc_hd__mux2_1 _09831_ (.A0(_05532_),
    .A1(\data_array.data0[12][56] ),
    .S(_03125_),
    .X(_01582_));
 sky130_fd_sc_hd__mux2_1 _09832_ (.A0(_05534_),
    .A1(\data_array.data0[12][57] ),
    .S(_03125_),
    .X(_01583_));
 sky130_fd_sc_hd__mux2_1 _09833_ (.A0(_05536_),
    .A1(\data_array.data0[12][58] ),
    .S(_03125_),
    .X(_01584_));
 sky130_fd_sc_hd__mux2_1 _09834_ (.A0(_05538_),
    .A1(\data_array.data0[12][59] ),
    .S(_03125_),
    .X(_01585_));
 sky130_fd_sc_hd__mux2_1 _09835_ (.A0(_05540_),
    .A1(\data_array.data0[12][60] ),
    .S(_03125_),
    .X(_01586_));
 sky130_fd_sc_hd__mux2_1 _09836_ (.A0(_05542_),
    .A1(\data_array.data0[12][61] ),
    .S(_03125_),
    .X(_01587_));
 sky130_fd_sc_hd__mux2_1 _09837_ (.A0(_05544_),
    .A1(\data_array.data0[12][62] ),
    .S(_03125_),
    .X(_01588_));
 sky130_fd_sc_hd__mux2_1 _09838_ (.A0(_05546_),
    .A1(\data_array.data0[12][63] ),
    .S(_03125_),
    .X(_01589_));
 sky130_fd_sc_hd__or2_2 _09839_ (.A(_05414_),
    .B(_05558_),
    .X(_03126_));
 sky130_fd_sc_hd__mux2_1 _09840_ (.A0(_05420_),
    .A1(\data_array.data0[13][0] ),
    .S(_03126_),
    .X(_01590_));
 sky130_fd_sc_hd__mux2_1 _09841_ (.A0(_05422_),
    .A1(\data_array.data0[13][1] ),
    .S(_03126_),
    .X(_01591_));
 sky130_fd_sc_hd__mux2_1 _09842_ (.A0(_05424_),
    .A1(\data_array.data0[13][2] ),
    .S(_03126_),
    .X(_01592_));
 sky130_fd_sc_hd__mux2_1 _09843_ (.A0(_05426_),
    .A1(\data_array.data0[13][3] ),
    .S(_03126_),
    .X(_01593_));
 sky130_fd_sc_hd__mux2_1 _09844_ (.A0(_05428_),
    .A1(\data_array.data0[13][4] ),
    .S(_03126_),
    .X(_01594_));
 sky130_fd_sc_hd__mux2_1 _09845_ (.A0(_05430_),
    .A1(\data_array.data0[13][5] ),
    .S(_03126_),
    .X(_01595_));
 sky130_fd_sc_hd__mux2_1 _09846_ (.A0(_05432_),
    .A1(\data_array.data0[13][6] ),
    .S(_03126_),
    .X(_01596_));
 sky130_fd_sc_hd__mux2_1 _09847_ (.A0(_05434_),
    .A1(\data_array.data0[13][7] ),
    .S(_03126_),
    .X(_01597_));
 sky130_fd_sc_hd__mux2_1 _09848_ (.A0(_05436_),
    .A1(\data_array.data0[13][8] ),
    .S(_03126_),
    .X(_01598_));
 sky130_fd_sc_hd__mux2_1 _09849_ (.A0(_05438_),
    .A1(\data_array.data0[13][9] ),
    .S(_03126_),
    .X(_01599_));
 sky130_fd_sc_hd__mux2_1 _09850_ (.A0(_05440_),
    .A1(\data_array.data0[13][10] ),
    .S(_03126_),
    .X(_01600_));
 sky130_fd_sc_hd__mux2_1 _09851_ (.A0(_05442_),
    .A1(\data_array.data0[13][11] ),
    .S(_03126_),
    .X(_01601_));
 sky130_fd_sc_hd__mux2_1 _09852_ (.A0(_05444_),
    .A1(\data_array.data0[13][12] ),
    .S(_03126_),
    .X(_01602_));
 sky130_fd_sc_hd__mux2_1 _09853_ (.A0(_05446_),
    .A1(\data_array.data0[13][13] ),
    .S(_03126_),
    .X(_01603_));
 sky130_fd_sc_hd__mux2_1 _09854_ (.A0(_05448_),
    .A1(\data_array.data0[13][14] ),
    .S(_03126_),
    .X(_01604_));
 sky130_fd_sc_hd__mux2_1 _09855_ (.A0(_05450_),
    .A1(\data_array.data0[13][15] ),
    .S(_03126_),
    .X(_01605_));
 sky130_fd_sc_hd__mux2_1 _09856_ (.A0(_05452_),
    .A1(\data_array.data0[13][16] ),
    .S(_03126_),
    .X(_01606_));
 sky130_fd_sc_hd__mux2_1 _09857_ (.A0(_05454_),
    .A1(\data_array.data0[13][17] ),
    .S(_03126_),
    .X(_01607_));
 sky130_fd_sc_hd__mux2_1 _09858_ (.A0(_05456_),
    .A1(\data_array.data0[13][18] ),
    .S(_03126_),
    .X(_01608_));
 sky130_fd_sc_hd__mux2_1 _09859_ (.A0(_05458_),
    .A1(\data_array.data0[13][19] ),
    .S(_03126_),
    .X(_01609_));
 sky130_fd_sc_hd__mux2_1 _09860_ (.A0(_05460_),
    .A1(\data_array.data0[13][20] ),
    .S(_03126_),
    .X(_01610_));
 sky130_fd_sc_hd__mux2_1 _09861_ (.A0(_05462_),
    .A1(\data_array.data0[13][21] ),
    .S(_03126_),
    .X(_01611_));
 sky130_fd_sc_hd__mux2_1 _09862_ (.A0(_05464_),
    .A1(\data_array.data0[13][22] ),
    .S(_03126_),
    .X(_01612_));
 sky130_fd_sc_hd__mux2_1 _09863_ (.A0(_05466_),
    .A1(\data_array.data0[13][23] ),
    .S(_03126_),
    .X(_01613_));
 sky130_fd_sc_hd__mux2_1 _09864_ (.A0(_05468_),
    .A1(\data_array.data0[13][24] ),
    .S(_03126_),
    .X(_01614_));
 sky130_fd_sc_hd__mux2_1 _09865_ (.A0(_05470_),
    .A1(\data_array.data0[13][25] ),
    .S(_03126_),
    .X(_01615_));
 sky130_fd_sc_hd__mux2_1 _09866_ (.A0(_05472_),
    .A1(\data_array.data0[13][26] ),
    .S(_03126_),
    .X(_01616_));
 sky130_fd_sc_hd__mux2_1 _09867_ (.A0(_05474_),
    .A1(\data_array.data0[13][27] ),
    .S(_03126_),
    .X(_01617_));
 sky130_fd_sc_hd__mux2_1 _09868_ (.A0(_05476_),
    .A1(\data_array.data0[13][28] ),
    .S(_03126_),
    .X(_01618_));
 sky130_fd_sc_hd__mux2_1 _09869_ (.A0(_05478_),
    .A1(\data_array.data0[13][29] ),
    .S(_03126_),
    .X(_01619_));
 sky130_fd_sc_hd__mux2_1 _09870_ (.A0(_05480_),
    .A1(\data_array.data0[13][30] ),
    .S(_03126_),
    .X(_01620_));
 sky130_fd_sc_hd__mux2_1 _09871_ (.A0(_05482_),
    .A1(\data_array.data0[13][31] ),
    .S(_03126_),
    .X(_01621_));
 sky130_fd_sc_hd__mux2_1 _09872_ (.A0(_05484_),
    .A1(\data_array.data0[13][32] ),
    .S(_03126_),
    .X(_01622_));
 sky130_fd_sc_hd__mux2_1 _09873_ (.A0(_05486_),
    .A1(\data_array.data0[13][33] ),
    .S(_03126_),
    .X(_01623_));
 sky130_fd_sc_hd__mux2_1 _09874_ (.A0(_05488_),
    .A1(\data_array.data0[13][34] ),
    .S(_03126_),
    .X(_01624_));
 sky130_fd_sc_hd__mux2_1 _09875_ (.A0(_05490_),
    .A1(\data_array.data0[13][35] ),
    .S(_03126_),
    .X(_01625_));
 sky130_fd_sc_hd__mux2_1 _09876_ (.A0(_05492_),
    .A1(\data_array.data0[13][36] ),
    .S(_03126_),
    .X(_01626_));
 sky130_fd_sc_hd__mux2_1 _09877_ (.A0(_05494_),
    .A1(\data_array.data0[13][37] ),
    .S(_03126_),
    .X(_01627_));
 sky130_fd_sc_hd__mux2_1 _09878_ (.A0(_05496_),
    .A1(\data_array.data0[13][38] ),
    .S(_03126_),
    .X(_01628_));
 sky130_fd_sc_hd__mux2_1 _09879_ (.A0(_05498_),
    .A1(\data_array.data0[13][39] ),
    .S(_03126_),
    .X(_01629_));
 sky130_fd_sc_hd__mux2_1 _09880_ (.A0(_05500_),
    .A1(\data_array.data0[13][40] ),
    .S(_03126_),
    .X(_01630_));
 sky130_fd_sc_hd__mux2_1 _09881_ (.A0(_05502_),
    .A1(\data_array.data0[13][41] ),
    .S(_03126_),
    .X(_01631_));
 sky130_fd_sc_hd__mux2_1 _09882_ (.A0(_05504_),
    .A1(\data_array.data0[13][42] ),
    .S(_03126_),
    .X(_01632_));
 sky130_fd_sc_hd__mux2_1 _09883_ (.A0(_05506_),
    .A1(\data_array.data0[13][43] ),
    .S(_03126_),
    .X(_01633_));
 sky130_fd_sc_hd__mux2_1 _09884_ (.A0(_05508_),
    .A1(\data_array.data0[13][44] ),
    .S(_03126_),
    .X(_01634_));
 sky130_fd_sc_hd__mux2_1 _09885_ (.A0(_05510_),
    .A1(\data_array.data0[13][45] ),
    .S(_03126_),
    .X(_01635_));
 sky130_fd_sc_hd__mux2_1 _09886_ (.A0(_05512_),
    .A1(\data_array.data0[13][46] ),
    .S(_03126_),
    .X(_01636_));
 sky130_fd_sc_hd__mux2_1 _09887_ (.A0(_05514_),
    .A1(\data_array.data0[13][47] ),
    .S(_03126_),
    .X(_01637_));
 sky130_fd_sc_hd__mux2_1 _09888_ (.A0(_05516_),
    .A1(\data_array.data0[13][48] ),
    .S(_03126_),
    .X(_01638_));
 sky130_fd_sc_hd__mux2_1 _09889_ (.A0(_05518_),
    .A1(\data_array.data0[13][49] ),
    .S(_03126_),
    .X(_01639_));
 sky130_fd_sc_hd__mux2_1 _09890_ (.A0(_05520_),
    .A1(\data_array.data0[13][50] ),
    .S(_03126_),
    .X(_01640_));
 sky130_fd_sc_hd__mux2_1 _09891_ (.A0(_05522_),
    .A1(\data_array.data0[13][51] ),
    .S(_03126_),
    .X(_01641_));
 sky130_fd_sc_hd__mux2_1 _09892_ (.A0(_05524_),
    .A1(\data_array.data0[13][52] ),
    .S(_03126_),
    .X(_01642_));
 sky130_fd_sc_hd__mux2_1 _09893_ (.A0(_05526_),
    .A1(\data_array.data0[13][53] ),
    .S(_03126_),
    .X(_01643_));
 sky130_fd_sc_hd__mux2_1 _09894_ (.A0(_05528_),
    .A1(\data_array.data0[13][54] ),
    .S(_03126_),
    .X(_01644_));
 sky130_fd_sc_hd__mux2_1 _09895_ (.A0(_05530_),
    .A1(\data_array.data0[13][55] ),
    .S(_03126_),
    .X(_01645_));
 sky130_fd_sc_hd__mux2_1 _09896_ (.A0(_05532_),
    .A1(\data_array.data0[13][56] ),
    .S(_03126_),
    .X(_01646_));
 sky130_fd_sc_hd__mux2_1 _09897_ (.A0(_05534_),
    .A1(\data_array.data0[13][57] ),
    .S(_03126_),
    .X(_01647_));
 sky130_fd_sc_hd__mux2_1 _09898_ (.A0(_05536_),
    .A1(\data_array.data0[13][58] ),
    .S(_03126_),
    .X(_01648_));
 sky130_fd_sc_hd__mux2_1 _09899_ (.A0(_05538_),
    .A1(\data_array.data0[13][59] ),
    .S(_03126_),
    .X(_01649_));
 sky130_fd_sc_hd__mux2_1 _09900_ (.A0(_05540_),
    .A1(\data_array.data0[13][60] ),
    .S(_03126_),
    .X(_01650_));
 sky130_fd_sc_hd__mux2_1 _09901_ (.A0(_05542_),
    .A1(\data_array.data0[13][61] ),
    .S(_03126_),
    .X(_01651_));
 sky130_fd_sc_hd__mux2_1 _09902_ (.A0(_05544_),
    .A1(\data_array.data0[13][62] ),
    .S(_03126_),
    .X(_01652_));
 sky130_fd_sc_hd__mux2_1 _09903_ (.A0(_05546_),
    .A1(\data_array.data0[13][63] ),
    .S(_03126_),
    .X(_01653_));
 sky130_fd_sc_hd__mux2_1 _09904_ (.A0(_05365_),
    .A1(\tag_array.tag0[4][0] ),
    .S(_05582_),
    .X(_01654_));
 sky130_fd_sc_hd__mux2_1 _09905_ (.A0(_05367_),
    .A1(\tag_array.tag0[4][1] ),
    .S(_05582_),
    .X(_01655_));
 sky130_fd_sc_hd__mux2_1 _09906_ (.A0(_05369_),
    .A1(\tag_array.tag0[4][2] ),
    .S(_05582_),
    .X(_01656_));
 sky130_fd_sc_hd__mux2_1 _09907_ (.A0(_05371_),
    .A1(\tag_array.tag0[4][3] ),
    .S(_05582_),
    .X(_01657_));
 sky130_fd_sc_hd__mux2_1 _09908_ (.A0(_05373_),
    .A1(\tag_array.tag0[4][4] ),
    .S(_05582_),
    .X(_01658_));
 sky130_fd_sc_hd__mux2_1 _09909_ (.A0(_05375_),
    .A1(\tag_array.tag0[4][5] ),
    .S(_05582_),
    .X(_01659_));
 sky130_fd_sc_hd__mux2_1 _09910_ (.A0(_05377_),
    .A1(\tag_array.tag0[4][6] ),
    .S(_05582_),
    .X(_01660_));
 sky130_fd_sc_hd__mux2_1 _09911_ (.A0(_05379_),
    .A1(\tag_array.tag0[4][7] ),
    .S(_05582_),
    .X(_01661_));
 sky130_fd_sc_hd__mux2_1 _09912_ (.A0(_05381_),
    .A1(\tag_array.tag0[4][8] ),
    .S(_05582_),
    .X(_01662_));
 sky130_fd_sc_hd__mux2_1 _09913_ (.A0(_05383_),
    .A1(\tag_array.tag0[4][9] ),
    .S(_05582_),
    .X(_01663_));
 sky130_fd_sc_hd__mux2_1 _09914_ (.A0(_05385_),
    .A1(\tag_array.tag0[4][10] ),
    .S(_05582_),
    .X(_01664_));
 sky130_fd_sc_hd__mux2_1 _09915_ (.A0(_05387_),
    .A1(\tag_array.tag0[4][11] ),
    .S(_05582_),
    .X(_01665_));
 sky130_fd_sc_hd__mux2_1 _09916_ (.A0(_05389_),
    .A1(\tag_array.tag0[4][12] ),
    .S(_05582_),
    .X(_01666_));
 sky130_fd_sc_hd__mux2_1 _09917_ (.A0(_05391_),
    .A1(\tag_array.tag0[4][13] ),
    .S(_05582_),
    .X(_01667_));
 sky130_fd_sc_hd__mux2_1 _09918_ (.A0(_05393_),
    .A1(\tag_array.tag0[4][14] ),
    .S(_05582_),
    .X(_01668_));
 sky130_fd_sc_hd__mux2_1 _09919_ (.A0(_05395_),
    .A1(\tag_array.tag0[4][15] ),
    .S(_05582_),
    .X(_01669_));
 sky130_fd_sc_hd__mux2_1 _09920_ (.A0(_05397_),
    .A1(\tag_array.tag0[4][16] ),
    .S(_05582_),
    .X(_01670_));
 sky130_fd_sc_hd__mux2_1 _09921_ (.A0(_05399_),
    .A1(\tag_array.tag0[4][17] ),
    .S(_05582_),
    .X(_01671_));
 sky130_fd_sc_hd__mux2_1 _09922_ (.A0(_05401_),
    .A1(\tag_array.tag0[4][18] ),
    .S(_05582_),
    .X(_01672_));
 sky130_fd_sc_hd__mux2_1 _09923_ (.A0(_05403_),
    .A1(\tag_array.tag0[4][19] ),
    .S(_05582_),
    .X(_01673_));
 sky130_fd_sc_hd__mux2_1 _09924_ (.A0(_05405_),
    .A1(\tag_array.tag0[4][20] ),
    .S(_05582_),
    .X(_01674_));
 sky130_fd_sc_hd__mux2_1 _09925_ (.A0(_05407_),
    .A1(\tag_array.tag0[4][21] ),
    .S(_05582_),
    .X(_01675_));
 sky130_fd_sc_hd__mux2_1 _09926_ (.A0(_05409_),
    .A1(\tag_array.tag0[4][22] ),
    .S(_05582_),
    .X(_01676_));
 sky130_fd_sc_hd__mux2_1 _09927_ (.A0(_05411_),
    .A1(\tag_array.tag0[4][23] ),
    .S(_05582_),
    .X(_01677_));
 sky130_fd_sc_hd__mux2_1 _09928_ (.A0(_05413_),
    .A1(\tag_array.tag0[4][24] ),
    .S(_05582_),
    .X(_01678_));
 sky130_fd_sc_hd__nand2_2 _09929_ (.A(_05415_),
    .B(_05583_),
    .Y(_03127_));
 sky130_fd_sc_hd__mux2_1 _09930_ (.A0(_05420_),
    .A1(\data_array.data0[3][0] ),
    .S(_03127_),
    .X(_01679_));
 sky130_fd_sc_hd__mux2_1 _09931_ (.A0(_05422_),
    .A1(\data_array.data0[3][1] ),
    .S(_03127_),
    .X(_01680_));
 sky130_fd_sc_hd__mux2_1 _09932_ (.A0(_05424_),
    .A1(\data_array.data0[3][2] ),
    .S(_03127_),
    .X(_01681_));
 sky130_fd_sc_hd__mux2_1 _09933_ (.A0(_05426_),
    .A1(\data_array.data0[3][3] ),
    .S(_03127_),
    .X(_01682_));
 sky130_fd_sc_hd__mux2_1 _09934_ (.A0(_05428_),
    .A1(\data_array.data0[3][4] ),
    .S(_03127_),
    .X(_01683_));
 sky130_fd_sc_hd__mux2_1 _09935_ (.A0(_05430_),
    .A1(\data_array.data0[3][5] ),
    .S(_03127_),
    .X(_01684_));
 sky130_fd_sc_hd__mux2_1 _09936_ (.A0(_05432_),
    .A1(\data_array.data0[3][6] ),
    .S(_03127_),
    .X(_01685_));
 sky130_fd_sc_hd__mux2_1 _09937_ (.A0(_05434_),
    .A1(\data_array.data0[3][7] ),
    .S(_03127_),
    .X(_01686_));
 sky130_fd_sc_hd__mux2_1 _09938_ (.A0(_05436_),
    .A1(\data_array.data0[3][8] ),
    .S(_03127_),
    .X(_01687_));
 sky130_fd_sc_hd__mux2_1 _09939_ (.A0(_05438_),
    .A1(\data_array.data0[3][9] ),
    .S(_03127_),
    .X(_01688_));
 sky130_fd_sc_hd__mux2_1 _09940_ (.A0(_05440_),
    .A1(\data_array.data0[3][10] ),
    .S(_03127_),
    .X(_01689_));
 sky130_fd_sc_hd__mux2_1 _09941_ (.A0(_05442_),
    .A1(\data_array.data0[3][11] ),
    .S(_03127_),
    .X(_01690_));
 sky130_fd_sc_hd__mux2_1 _09942_ (.A0(_05444_),
    .A1(\data_array.data0[3][12] ),
    .S(_03127_),
    .X(_01691_));
 sky130_fd_sc_hd__mux2_1 _09943_ (.A0(_05446_),
    .A1(\data_array.data0[3][13] ),
    .S(_03127_),
    .X(_01692_));
 sky130_fd_sc_hd__mux2_1 _09944_ (.A0(_05448_),
    .A1(\data_array.data0[3][14] ),
    .S(_03127_),
    .X(_01693_));
 sky130_fd_sc_hd__mux2_1 _09945_ (.A0(_05450_),
    .A1(\data_array.data0[3][15] ),
    .S(_03127_),
    .X(_01694_));
 sky130_fd_sc_hd__mux2_1 _09946_ (.A0(_05452_),
    .A1(\data_array.data0[3][16] ),
    .S(_03127_),
    .X(_01695_));
 sky130_fd_sc_hd__mux2_1 _09947_ (.A0(_05454_),
    .A1(\data_array.data0[3][17] ),
    .S(_03127_),
    .X(_01696_));
 sky130_fd_sc_hd__mux2_1 _09948_ (.A0(_05456_),
    .A1(\data_array.data0[3][18] ),
    .S(_03127_),
    .X(_01697_));
 sky130_fd_sc_hd__mux2_1 _09949_ (.A0(_05458_),
    .A1(\data_array.data0[3][19] ),
    .S(_03127_),
    .X(_01698_));
 sky130_fd_sc_hd__mux2_1 _09950_ (.A0(_05460_),
    .A1(\data_array.data0[3][20] ),
    .S(_03127_),
    .X(_01699_));
 sky130_fd_sc_hd__mux2_1 _09951_ (.A0(_05462_),
    .A1(\data_array.data0[3][21] ),
    .S(_03127_),
    .X(_01700_));
 sky130_fd_sc_hd__mux2_1 _09952_ (.A0(_05464_),
    .A1(\data_array.data0[3][22] ),
    .S(_03127_),
    .X(_01701_));
 sky130_fd_sc_hd__mux2_1 _09953_ (.A0(_05466_),
    .A1(\data_array.data0[3][23] ),
    .S(_03127_),
    .X(_01702_));
 sky130_fd_sc_hd__mux2_1 _09954_ (.A0(_05468_),
    .A1(\data_array.data0[3][24] ),
    .S(_03127_),
    .X(_01703_));
 sky130_fd_sc_hd__mux2_1 _09955_ (.A0(_05470_),
    .A1(\data_array.data0[3][25] ),
    .S(_03127_),
    .X(_01704_));
 sky130_fd_sc_hd__mux2_1 _09956_ (.A0(_05472_),
    .A1(\data_array.data0[3][26] ),
    .S(_03127_),
    .X(_01705_));
 sky130_fd_sc_hd__mux2_1 _09957_ (.A0(_05474_),
    .A1(\data_array.data0[3][27] ),
    .S(_03127_),
    .X(_01706_));
 sky130_fd_sc_hd__mux2_1 _09958_ (.A0(_05476_),
    .A1(\data_array.data0[3][28] ),
    .S(_03127_),
    .X(_01707_));
 sky130_fd_sc_hd__mux2_1 _09959_ (.A0(_05478_),
    .A1(\data_array.data0[3][29] ),
    .S(_03127_),
    .X(_01708_));
 sky130_fd_sc_hd__mux2_1 _09960_ (.A0(_05480_),
    .A1(\data_array.data0[3][30] ),
    .S(_03127_),
    .X(_01709_));
 sky130_fd_sc_hd__mux2_1 _09961_ (.A0(_05482_),
    .A1(\data_array.data0[3][31] ),
    .S(_03127_),
    .X(_01710_));
 sky130_fd_sc_hd__mux2_1 _09962_ (.A0(_05484_),
    .A1(\data_array.data0[3][32] ),
    .S(_03127_),
    .X(_01711_));
 sky130_fd_sc_hd__mux2_1 _09963_ (.A0(_05486_),
    .A1(\data_array.data0[3][33] ),
    .S(_03127_),
    .X(_01712_));
 sky130_fd_sc_hd__mux2_1 _09964_ (.A0(_05488_),
    .A1(\data_array.data0[3][34] ),
    .S(_03127_),
    .X(_01713_));
 sky130_fd_sc_hd__mux2_1 _09965_ (.A0(_05490_),
    .A1(\data_array.data0[3][35] ),
    .S(_03127_),
    .X(_01714_));
 sky130_fd_sc_hd__mux2_1 _09966_ (.A0(_05492_),
    .A1(\data_array.data0[3][36] ),
    .S(_03127_),
    .X(_01715_));
 sky130_fd_sc_hd__mux2_1 _09967_ (.A0(_05494_),
    .A1(\data_array.data0[3][37] ),
    .S(_03127_),
    .X(_01716_));
 sky130_fd_sc_hd__mux2_1 _09968_ (.A0(_05496_),
    .A1(\data_array.data0[3][38] ),
    .S(_03127_),
    .X(_01717_));
 sky130_fd_sc_hd__mux2_1 _09969_ (.A0(_05498_),
    .A1(\data_array.data0[3][39] ),
    .S(_03127_),
    .X(_01718_));
 sky130_fd_sc_hd__mux2_1 _09970_ (.A0(_05500_),
    .A1(\data_array.data0[3][40] ),
    .S(_03127_),
    .X(_01719_));
 sky130_fd_sc_hd__mux2_1 _09971_ (.A0(_05502_),
    .A1(\data_array.data0[3][41] ),
    .S(_03127_),
    .X(_01720_));
 sky130_fd_sc_hd__mux2_1 _09972_ (.A0(_05504_),
    .A1(\data_array.data0[3][42] ),
    .S(_03127_),
    .X(_01721_));
 sky130_fd_sc_hd__mux2_1 _09973_ (.A0(_05506_),
    .A1(\data_array.data0[3][43] ),
    .S(_03127_),
    .X(_01722_));
 sky130_fd_sc_hd__mux2_1 _09974_ (.A0(_05508_),
    .A1(\data_array.data0[3][44] ),
    .S(_03127_),
    .X(_01723_));
 sky130_fd_sc_hd__mux2_1 _09975_ (.A0(_05510_),
    .A1(\data_array.data0[3][45] ),
    .S(_03127_),
    .X(_01724_));
 sky130_fd_sc_hd__mux2_1 _09976_ (.A0(_05512_),
    .A1(\data_array.data0[3][46] ),
    .S(_03127_),
    .X(_01725_));
 sky130_fd_sc_hd__mux2_1 _09977_ (.A0(_05514_),
    .A1(\data_array.data0[3][47] ),
    .S(_03127_),
    .X(_01726_));
 sky130_fd_sc_hd__mux2_1 _09978_ (.A0(_05516_),
    .A1(\data_array.data0[3][48] ),
    .S(_03127_),
    .X(_01727_));
 sky130_fd_sc_hd__mux2_1 _09979_ (.A0(_05518_),
    .A1(\data_array.data0[3][49] ),
    .S(_03127_),
    .X(_01728_));
 sky130_fd_sc_hd__mux2_1 _09980_ (.A0(_05520_),
    .A1(\data_array.data0[3][50] ),
    .S(_03127_),
    .X(_01729_));
 sky130_fd_sc_hd__mux2_1 _09981_ (.A0(_05522_),
    .A1(\data_array.data0[3][51] ),
    .S(_03127_),
    .X(_01730_));
 sky130_fd_sc_hd__mux2_1 _09982_ (.A0(_05524_),
    .A1(\data_array.data0[3][52] ),
    .S(_03127_),
    .X(_01731_));
 sky130_fd_sc_hd__mux2_1 _09983_ (.A0(_05526_),
    .A1(\data_array.data0[3][53] ),
    .S(_03127_),
    .X(_01732_));
 sky130_fd_sc_hd__mux2_1 _09984_ (.A0(_05528_),
    .A1(\data_array.data0[3][54] ),
    .S(_03127_),
    .X(_01733_));
 sky130_fd_sc_hd__mux2_1 _09985_ (.A0(_05530_),
    .A1(\data_array.data0[3][55] ),
    .S(_03127_),
    .X(_01734_));
 sky130_fd_sc_hd__mux2_1 _09986_ (.A0(_05532_),
    .A1(\data_array.data0[3][56] ),
    .S(_03127_),
    .X(_01735_));
 sky130_fd_sc_hd__mux2_1 _09987_ (.A0(_05534_),
    .A1(\data_array.data0[3][57] ),
    .S(_03127_),
    .X(_01736_));
 sky130_fd_sc_hd__mux2_1 _09988_ (.A0(_05536_),
    .A1(\data_array.data0[3][58] ),
    .S(_03127_),
    .X(_01737_));
 sky130_fd_sc_hd__mux2_1 _09989_ (.A0(_05538_),
    .A1(\data_array.data0[3][59] ),
    .S(_03127_),
    .X(_01738_));
 sky130_fd_sc_hd__mux2_1 _09990_ (.A0(_05540_),
    .A1(\data_array.data0[3][60] ),
    .S(_03127_),
    .X(_01739_));
 sky130_fd_sc_hd__mux2_1 _09991_ (.A0(_05542_),
    .A1(\data_array.data0[3][61] ),
    .S(_03127_),
    .X(_01740_));
 sky130_fd_sc_hd__mux2_1 _09992_ (.A0(_05544_),
    .A1(\data_array.data0[3][62] ),
    .S(_03127_),
    .X(_01741_));
 sky130_fd_sc_hd__mux2_1 _09993_ (.A0(_05546_),
    .A1(\data_array.data0[3][63] ),
    .S(_03127_),
    .X(_01742_));
 sky130_fd_sc_hd__mux2_1 _09994_ (.A0(_05420_),
    .A1(\data_array.data1[13][0] ),
    .S(_05593_),
    .X(_01743_));
 sky130_fd_sc_hd__mux2_1 _09995_ (.A0(_05422_),
    .A1(\data_array.data1[13][1] ),
    .S(_05593_),
    .X(_01744_));
 sky130_fd_sc_hd__mux2_1 _09996_ (.A0(_05424_),
    .A1(\data_array.data1[13][2] ),
    .S(_05593_),
    .X(_01745_));
 sky130_fd_sc_hd__mux2_1 _09997_ (.A0(_05426_),
    .A1(\data_array.data1[13][3] ),
    .S(_05593_),
    .X(_01746_));
 sky130_fd_sc_hd__mux2_1 _09998_ (.A0(_05428_),
    .A1(\data_array.data1[13][4] ),
    .S(_05593_),
    .X(_01747_));
 sky130_fd_sc_hd__mux2_1 _09999_ (.A0(_05430_),
    .A1(\data_array.data1[13][5] ),
    .S(_05593_),
    .X(_01748_));
 sky130_fd_sc_hd__mux2_1 _10000_ (.A0(_05432_),
    .A1(\data_array.data1[13][6] ),
    .S(_05593_),
    .X(_01749_));
 sky130_fd_sc_hd__mux2_1 _10001_ (.A0(_05434_),
    .A1(\data_array.data1[13][7] ),
    .S(_05593_),
    .X(_01750_));
 sky130_fd_sc_hd__mux2_1 _10002_ (.A0(_05436_),
    .A1(\data_array.data1[13][8] ),
    .S(_05593_),
    .X(_01751_));
 sky130_fd_sc_hd__mux2_1 _10003_ (.A0(_05438_),
    .A1(\data_array.data1[13][9] ),
    .S(_05593_),
    .X(_01752_));
 sky130_fd_sc_hd__mux2_1 _10004_ (.A0(_05440_),
    .A1(\data_array.data1[13][10] ),
    .S(_05593_),
    .X(_01753_));
 sky130_fd_sc_hd__mux2_1 _10005_ (.A0(_05442_),
    .A1(\data_array.data1[13][11] ),
    .S(_05593_),
    .X(_01754_));
 sky130_fd_sc_hd__mux2_1 _10006_ (.A0(_05444_),
    .A1(\data_array.data1[13][12] ),
    .S(_05593_),
    .X(_01755_));
 sky130_fd_sc_hd__mux2_1 _10007_ (.A0(_05446_),
    .A1(\data_array.data1[13][13] ),
    .S(_05593_),
    .X(_01756_));
 sky130_fd_sc_hd__mux2_1 _10008_ (.A0(_05448_),
    .A1(\data_array.data1[13][14] ),
    .S(_05593_),
    .X(_01757_));
 sky130_fd_sc_hd__mux2_1 _10009_ (.A0(_05450_),
    .A1(\data_array.data1[13][15] ),
    .S(_05593_),
    .X(_01758_));
 sky130_fd_sc_hd__mux2_1 _10010_ (.A0(_05452_),
    .A1(\data_array.data1[13][16] ),
    .S(_05593_),
    .X(_01759_));
 sky130_fd_sc_hd__mux2_1 _10011_ (.A0(_05454_),
    .A1(\data_array.data1[13][17] ),
    .S(_05593_),
    .X(_01760_));
 sky130_fd_sc_hd__mux2_1 _10012_ (.A0(_05456_),
    .A1(\data_array.data1[13][18] ),
    .S(_05593_),
    .X(_01761_));
 sky130_fd_sc_hd__mux2_1 _10013_ (.A0(_05458_),
    .A1(\data_array.data1[13][19] ),
    .S(_05593_),
    .X(_01762_));
 sky130_fd_sc_hd__mux2_1 _10014_ (.A0(_05460_),
    .A1(\data_array.data1[13][20] ),
    .S(_05593_),
    .X(_01763_));
 sky130_fd_sc_hd__mux2_1 _10015_ (.A0(_05462_),
    .A1(\data_array.data1[13][21] ),
    .S(_05593_),
    .X(_01764_));
 sky130_fd_sc_hd__mux2_1 _10016_ (.A0(_05464_),
    .A1(\data_array.data1[13][22] ),
    .S(_05593_),
    .X(_01765_));
 sky130_fd_sc_hd__mux2_1 _10017_ (.A0(_05466_),
    .A1(\data_array.data1[13][23] ),
    .S(_05593_),
    .X(_01766_));
 sky130_fd_sc_hd__mux2_1 _10018_ (.A0(_05468_),
    .A1(\data_array.data1[13][24] ),
    .S(_05593_),
    .X(_01767_));
 sky130_fd_sc_hd__mux2_1 _10019_ (.A0(_05470_),
    .A1(\data_array.data1[13][25] ),
    .S(_05593_),
    .X(_01768_));
 sky130_fd_sc_hd__mux2_1 _10020_ (.A0(_05472_),
    .A1(\data_array.data1[13][26] ),
    .S(_05593_),
    .X(_01769_));
 sky130_fd_sc_hd__mux2_1 _10021_ (.A0(_05474_),
    .A1(\data_array.data1[13][27] ),
    .S(_05593_),
    .X(_01770_));
 sky130_fd_sc_hd__mux2_1 _10022_ (.A0(_05476_),
    .A1(\data_array.data1[13][28] ),
    .S(_05593_),
    .X(_01771_));
 sky130_fd_sc_hd__mux2_1 _10023_ (.A0(_05478_),
    .A1(\data_array.data1[13][29] ),
    .S(_05593_),
    .X(_01772_));
 sky130_fd_sc_hd__mux2_1 _10024_ (.A0(_05480_),
    .A1(\data_array.data1[13][30] ),
    .S(_05593_),
    .X(_01773_));
 sky130_fd_sc_hd__mux2_1 _10025_ (.A0(_05482_),
    .A1(\data_array.data1[13][31] ),
    .S(_05593_),
    .X(_01774_));
 sky130_fd_sc_hd__mux2_1 _10026_ (.A0(_05484_),
    .A1(\data_array.data1[13][32] ),
    .S(_05593_),
    .X(_01775_));
 sky130_fd_sc_hd__mux2_1 _10027_ (.A0(_05486_),
    .A1(\data_array.data1[13][33] ),
    .S(_05593_),
    .X(_01776_));
 sky130_fd_sc_hd__mux2_1 _10028_ (.A0(_05488_),
    .A1(\data_array.data1[13][34] ),
    .S(_05593_),
    .X(_01777_));
 sky130_fd_sc_hd__mux2_1 _10029_ (.A0(_05490_),
    .A1(\data_array.data1[13][35] ),
    .S(_05593_),
    .X(_01778_));
 sky130_fd_sc_hd__mux2_1 _10030_ (.A0(_05492_),
    .A1(\data_array.data1[13][36] ),
    .S(_05593_),
    .X(_01779_));
 sky130_fd_sc_hd__mux2_1 _10031_ (.A0(_05494_),
    .A1(\data_array.data1[13][37] ),
    .S(_05593_),
    .X(_01780_));
 sky130_fd_sc_hd__mux2_1 _10032_ (.A0(_05496_),
    .A1(\data_array.data1[13][38] ),
    .S(_05593_),
    .X(_01781_));
 sky130_fd_sc_hd__mux2_1 _10033_ (.A0(_05498_),
    .A1(\data_array.data1[13][39] ),
    .S(_05593_),
    .X(_01782_));
 sky130_fd_sc_hd__mux2_1 _10034_ (.A0(_05500_),
    .A1(\data_array.data1[13][40] ),
    .S(_05593_),
    .X(_01783_));
 sky130_fd_sc_hd__mux2_1 _10035_ (.A0(_05502_),
    .A1(\data_array.data1[13][41] ),
    .S(_05593_),
    .X(_01784_));
 sky130_fd_sc_hd__mux2_1 _10036_ (.A0(_05504_),
    .A1(\data_array.data1[13][42] ),
    .S(_05593_),
    .X(_01785_));
 sky130_fd_sc_hd__mux2_1 _10037_ (.A0(_05506_),
    .A1(\data_array.data1[13][43] ),
    .S(_05593_),
    .X(_01786_));
 sky130_fd_sc_hd__mux2_1 _10038_ (.A0(_05508_),
    .A1(\data_array.data1[13][44] ),
    .S(_05593_),
    .X(_01787_));
 sky130_fd_sc_hd__mux2_1 _10039_ (.A0(_05510_),
    .A1(\data_array.data1[13][45] ),
    .S(_05593_),
    .X(_01788_));
 sky130_fd_sc_hd__mux2_1 _10040_ (.A0(_05512_),
    .A1(\data_array.data1[13][46] ),
    .S(_05593_),
    .X(_01789_));
 sky130_fd_sc_hd__mux2_1 _10041_ (.A0(_05514_),
    .A1(\data_array.data1[13][47] ),
    .S(_05593_),
    .X(_01790_));
 sky130_fd_sc_hd__mux2_1 _10042_ (.A0(_05516_),
    .A1(\data_array.data1[13][48] ),
    .S(_05593_),
    .X(_01791_));
 sky130_fd_sc_hd__mux2_1 _10043_ (.A0(_05518_),
    .A1(\data_array.data1[13][49] ),
    .S(_05593_),
    .X(_01792_));
 sky130_fd_sc_hd__mux2_1 _10044_ (.A0(_05520_),
    .A1(\data_array.data1[13][50] ),
    .S(_05593_),
    .X(_01793_));
 sky130_fd_sc_hd__mux2_1 _10045_ (.A0(_05522_),
    .A1(\data_array.data1[13][51] ),
    .S(_05593_),
    .X(_01794_));
 sky130_fd_sc_hd__mux2_1 _10046_ (.A0(_05524_),
    .A1(\data_array.data1[13][52] ),
    .S(_05593_),
    .X(_01795_));
 sky130_fd_sc_hd__mux2_1 _10047_ (.A0(_05526_),
    .A1(\data_array.data1[13][53] ),
    .S(_05593_),
    .X(_01796_));
 sky130_fd_sc_hd__mux2_1 _10048_ (.A0(_05528_),
    .A1(\data_array.data1[13][54] ),
    .S(_05593_),
    .X(_01797_));
 sky130_fd_sc_hd__mux2_1 _10049_ (.A0(_05530_),
    .A1(\data_array.data1[13][55] ),
    .S(_05593_),
    .X(_01798_));
 sky130_fd_sc_hd__mux2_1 _10050_ (.A0(_05532_),
    .A1(\data_array.data1[13][56] ),
    .S(_05593_),
    .X(_01799_));
 sky130_fd_sc_hd__mux2_1 _10051_ (.A0(_05534_),
    .A1(\data_array.data1[13][57] ),
    .S(_05593_),
    .X(_01800_));
 sky130_fd_sc_hd__mux2_1 _10052_ (.A0(_05536_),
    .A1(\data_array.data1[13][58] ),
    .S(_05593_),
    .X(_01801_));
 sky130_fd_sc_hd__mux2_1 _10053_ (.A0(_05538_),
    .A1(\data_array.data1[13][59] ),
    .S(_05593_),
    .X(_01802_));
 sky130_fd_sc_hd__mux2_1 _10054_ (.A0(_05540_),
    .A1(\data_array.data1[13][60] ),
    .S(_05593_),
    .X(_01803_));
 sky130_fd_sc_hd__mux2_1 _10055_ (.A0(_05542_),
    .A1(\data_array.data1[13][61] ),
    .S(_05593_),
    .X(_01804_));
 sky130_fd_sc_hd__mux2_1 _10056_ (.A0(_05544_),
    .A1(\data_array.data1[13][62] ),
    .S(_05593_),
    .X(_01805_));
 sky130_fd_sc_hd__mux2_1 _10057_ (.A0(_05546_),
    .A1(\data_array.data1[13][63] ),
    .S(_05593_),
    .X(_01806_));
 sky130_fd_sc_hd__mux2_1 _10058_ (.A0(_05365_),
    .A1(\tag_array.tag0[3][0] ),
    .S(_05585_),
    .X(_01807_));
 sky130_fd_sc_hd__mux2_1 _10059_ (.A0(_05367_),
    .A1(\tag_array.tag0[3][1] ),
    .S(_05585_),
    .X(_01808_));
 sky130_fd_sc_hd__mux2_1 _10060_ (.A0(_05369_),
    .A1(\tag_array.tag0[3][2] ),
    .S(_05585_),
    .X(_01809_));
 sky130_fd_sc_hd__mux2_1 _10061_ (.A0(_05371_),
    .A1(\tag_array.tag0[3][3] ),
    .S(_05585_),
    .X(_01810_));
 sky130_fd_sc_hd__mux2_1 _10062_ (.A0(_05373_),
    .A1(\tag_array.tag0[3][4] ),
    .S(_05585_),
    .X(_01811_));
 sky130_fd_sc_hd__mux2_1 _10063_ (.A0(_05375_),
    .A1(\tag_array.tag0[3][5] ),
    .S(_05585_),
    .X(_01812_));
 sky130_fd_sc_hd__mux2_1 _10064_ (.A0(_05377_),
    .A1(\tag_array.tag0[3][6] ),
    .S(_05585_),
    .X(_01813_));
 sky130_fd_sc_hd__mux2_1 _10065_ (.A0(_05379_),
    .A1(\tag_array.tag0[3][7] ),
    .S(_05585_),
    .X(_01814_));
 sky130_fd_sc_hd__mux2_1 _10066_ (.A0(_05381_),
    .A1(\tag_array.tag0[3][8] ),
    .S(_05585_),
    .X(_01815_));
 sky130_fd_sc_hd__mux2_1 _10067_ (.A0(_05383_),
    .A1(\tag_array.tag0[3][9] ),
    .S(_05585_),
    .X(_01816_));
 sky130_fd_sc_hd__mux2_1 _10068_ (.A0(_05385_),
    .A1(\tag_array.tag0[3][10] ),
    .S(_05585_),
    .X(_01817_));
 sky130_fd_sc_hd__mux2_1 _10069_ (.A0(_05387_),
    .A1(\tag_array.tag0[3][11] ),
    .S(_05585_),
    .X(_01818_));
 sky130_fd_sc_hd__mux2_1 _10070_ (.A0(_05389_),
    .A1(\tag_array.tag0[3][12] ),
    .S(_05585_),
    .X(_01819_));
 sky130_fd_sc_hd__mux2_1 _10071_ (.A0(_05391_),
    .A1(\tag_array.tag0[3][13] ),
    .S(_05585_),
    .X(_01820_));
 sky130_fd_sc_hd__mux2_1 _10072_ (.A0(_05393_),
    .A1(\tag_array.tag0[3][14] ),
    .S(_05585_),
    .X(_01821_));
 sky130_fd_sc_hd__mux2_1 _10073_ (.A0(_05395_),
    .A1(\tag_array.tag0[3][15] ),
    .S(_05585_),
    .X(_01822_));
 sky130_fd_sc_hd__mux2_1 _10074_ (.A0(_05397_),
    .A1(\tag_array.tag0[3][16] ),
    .S(_05585_),
    .X(_01823_));
 sky130_fd_sc_hd__mux2_1 _10075_ (.A0(_05399_),
    .A1(\tag_array.tag0[3][17] ),
    .S(_05585_),
    .X(_01824_));
 sky130_fd_sc_hd__mux2_1 _10076_ (.A0(_05401_),
    .A1(\tag_array.tag0[3][18] ),
    .S(_05585_),
    .X(_01825_));
 sky130_fd_sc_hd__mux2_1 _10077_ (.A0(_05403_),
    .A1(\tag_array.tag0[3][19] ),
    .S(_05585_),
    .X(_01826_));
 sky130_fd_sc_hd__mux2_1 _10078_ (.A0(_05405_),
    .A1(\tag_array.tag0[3][20] ),
    .S(_05585_),
    .X(_01827_));
 sky130_fd_sc_hd__mux2_1 _10079_ (.A0(_05407_),
    .A1(\tag_array.tag0[3][21] ),
    .S(_05585_),
    .X(_01828_));
 sky130_fd_sc_hd__mux2_1 _10080_ (.A0(_05409_),
    .A1(\tag_array.tag0[3][22] ),
    .S(_05585_),
    .X(_01829_));
 sky130_fd_sc_hd__mux2_1 _10081_ (.A0(_05411_),
    .A1(\tag_array.tag0[3][23] ),
    .S(_05585_),
    .X(_01830_));
 sky130_fd_sc_hd__mux2_1 _10082_ (.A0(_05413_),
    .A1(\tag_array.tag0[3][24] ),
    .S(_05585_),
    .X(_01831_));
 sky130_fd_sc_hd__mux2_1 _10083_ (.A0(\tag_array.tag1[8][0] ),
    .A1(_05365_),
    .S(_05557_),
    .X(_01832_));
 sky130_fd_sc_hd__mux2_1 _10084_ (.A0(\tag_array.tag1[8][1] ),
    .A1(_05367_),
    .S(_05557_),
    .X(_01833_));
 sky130_fd_sc_hd__mux2_1 _10085_ (.A0(\tag_array.tag1[8][2] ),
    .A1(_05369_),
    .S(_05557_),
    .X(_01834_));
 sky130_fd_sc_hd__mux2_1 _10086_ (.A0(\tag_array.tag1[8][3] ),
    .A1(_05371_),
    .S(_05557_),
    .X(_01835_));
 sky130_fd_sc_hd__mux2_1 _10087_ (.A0(\tag_array.tag1[8][4] ),
    .A1(_05373_),
    .S(_05557_),
    .X(_01836_));
 sky130_fd_sc_hd__mux2_1 _10088_ (.A0(\tag_array.tag1[8][5] ),
    .A1(_05375_),
    .S(_05557_),
    .X(_01837_));
 sky130_fd_sc_hd__mux2_1 _10089_ (.A0(\tag_array.tag1[8][6] ),
    .A1(_05377_),
    .S(_05557_),
    .X(_01838_));
 sky130_fd_sc_hd__mux2_1 _10090_ (.A0(\tag_array.tag1[8][7] ),
    .A1(_05379_),
    .S(_05557_),
    .X(_01839_));
 sky130_fd_sc_hd__mux2_1 _10091_ (.A0(\tag_array.tag1[8][8] ),
    .A1(_05381_),
    .S(_05557_),
    .X(_01840_));
 sky130_fd_sc_hd__mux2_1 _10092_ (.A0(\tag_array.tag1[8][9] ),
    .A1(_05383_),
    .S(_05557_),
    .X(_01841_));
 sky130_fd_sc_hd__mux2_1 _10093_ (.A0(\tag_array.tag1[8][10] ),
    .A1(_05385_),
    .S(_05557_),
    .X(_01842_));
 sky130_fd_sc_hd__mux2_1 _10094_ (.A0(\tag_array.tag1[8][11] ),
    .A1(_05387_),
    .S(_05557_),
    .X(_01843_));
 sky130_fd_sc_hd__mux2_1 _10095_ (.A0(\tag_array.tag1[8][12] ),
    .A1(_05389_),
    .S(_05557_),
    .X(_01844_));
 sky130_fd_sc_hd__mux2_1 _10096_ (.A0(\tag_array.tag1[8][13] ),
    .A1(_05391_),
    .S(_05557_),
    .X(_01845_));
 sky130_fd_sc_hd__mux2_1 _10097_ (.A0(\tag_array.tag1[8][14] ),
    .A1(_05393_),
    .S(_05557_),
    .X(_01846_));
 sky130_fd_sc_hd__mux2_1 _10098_ (.A0(\tag_array.tag1[8][15] ),
    .A1(_05395_),
    .S(_05557_),
    .X(_01847_));
 sky130_fd_sc_hd__mux2_1 _10099_ (.A0(\tag_array.tag1[8][16] ),
    .A1(_05397_),
    .S(_05557_),
    .X(_01848_));
 sky130_fd_sc_hd__mux2_1 _10100_ (.A0(\tag_array.tag1[8][17] ),
    .A1(_05399_),
    .S(_05557_),
    .X(_01849_));
 sky130_fd_sc_hd__mux2_1 _10101_ (.A0(\tag_array.tag1[8][18] ),
    .A1(_05401_),
    .S(_05557_),
    .X(_01850_));
 sky130_fd_sc_hd__mux2_1 _10102_ (.A0(\tag_array.tag1[8][19] ),
    .A1(_05403_),
    .S(_05557_),
    .X(_01851_));
 sky130_fd_sc_hd__mux2_1 _10103_ (.A0(\tag_array.tag1[8][20] ),
    .A1(_05405_),
    .S(_05557_),
    .X(_01852_));
 sky130_fd_sc_hd__mux2_1 _10104_ (.A0(\tag_array.tag1[8][21] ),
    .A1(_05407_),
    .S(_05557_),
    .X(_01853_));
 sky130_fd_sc_hd__mux2_1 _10105_ (.A0(\tag_array.tag1[8][22] ),
    .A1(_05409_),
    .S(_05557_),
    .X(_01854_));
 sky130_fd_sc_hd__mux2_1 _10106_ (.A0(\tag_array.tag1[8][23] ),
    .A1(_05411_),
    .S(_05557_),
    .X(_01855_));
 sky130_fd_sc_hd__mux2_1 _10107_ (.A0(\tag_array.tag1[8][24] ),
    .A1(_05413_),
    .S(_05557_),
    .X(_01856_));
 sky130_fd_sc_hd__or2_2 _10108_ (.A(_05414_),
    .B(_05550_),
    .X(_03128_));
 sky130_fd_sc_hd__mux2_1 _10109_ (.A0(_05420_),
    .A1(\data_array.data0[11][0] ),
    .S(_03128_),
    .X(_01857_));
 sky130_fd_sc_hd__mux2_1 _10110_ (.A0(_05422_),
    .A1(\data_array.data0[11][1] ),
    .S(_03128_),
    .X(_01858_));
 sky130_fd_sc_hd__mux2_1 _10111_ (.A0(_05424_),
    .A1(\data_array.data0[11][2] ),
    .S(_03128_),
    .X(_01859_));
 sky130_fd_sc_hd__mux2_1 _10112_ (.A0(_05426_),
    .A1(\data_array.data0[11][3] ),
    .S(_03128_),
    .X(_01860_));
 sky130_fd_sc_hd__mux2_1 _10113_ (.A0(_05428_),
    .A1(\data_array.data0[11][4] ),
    .S(_03128_),
    .X(_01861_));
 sky130_fd_sc_hd__mux2_1 _10114_ (.A0(_05430_),
    .A1(\data_array.data0[11][5] ),
    .S(_03128_),
    .X(_01862_));
 sky130_fd_sc_hd__mux2_1 _10115_ (.A0(_05432_),
    .A1(\data_array.data0[11][6] ),
    .S(_03128_),
    .X(_01863_));
 sky130_fd_sc_hd__mux2_1 _10116_ (.A0(_05434_),
    .A1(\data_array.data0[11][7] ),
    .S(_03128_),
    .X(_01864_));
 sky130_fd_sc_hd__mux2_1 _10117_ (.A0(_05436_),
    .A1(\data_array.data0[11][8] ),
    .S(_03128_),
    .X(_01865_));
 sky130_fd_sc_hd__mux2_1 _10118_ (.A0(_05438_),
    .A1(\data_array.data0[11][9] ),
    .S(_03128_),
    .X(_01866_));
 sky130_fd_sc_hd__mux2_1 _10119_ (.A0(_05440_),
    .A1(\data_array.data0[11][10] ),
    .S(_03128_),
    .X(_01867_));
 sky130_fd_sc_hd__mux2_1 _10120_ (.A0(_05442_),
    .A1(\data_array.data0[11][11] ),
    .S(_03128_),
    .X(_01868_));
 sky130_fd_sc_hd__mux2_1 _10121_ (.A0(_05444_),
    .A1(\data_array.data0[11][12] ),
    .S(_03128_),
    .X(_01869_));
 sky130_fd_sc_hd__mux2_1 _10122_ (.A0(_05446_),
    .A1(\data_array.data0[11][13] ),
    .S(_03128_),
    .X(_01870_));
 sky130_fd_sc_hd__mux2_1 _10123_ (.A0(_05448_),
    .A1(\data_array.data0[11][14] ),
    .S(_03128_),
    .X(_01871_));
 sky130_fd_sc_hd__mux2_1 _10124_ (.A0(_05450_),
    .A1(\data_array.data0[11][15] ),
    .S(_03128_),
    .X(_01872_));
 sky130_fd_sc_hd__mux2_1 _10125_ (.A0(_05452_),
    .A1(\data_array.data0[11][16] ),
    .S(_03128_),
    .X(_01873_));
 sky130_fd_sc_hd__mux2_1 _10126_ (.A0(_05454_),
    .A1(\data_array.data0[11][17] ),
    .S(_03128_),
    .X(_01874_));
 sky130_fd_sc_hd__mux2_1 _10127_ (.A0(_05456_),
    .A1(\data_array.data0[11][18] ),
    .S(_03128_),
    .X(_01875_));
 sky130_fd_sc_hd__mux2_1 _10128_ (.A0(_05458_),
    .A1(\data_array.data0[11][19] ),
    .S(_03128_),
    .X(_01876_));
 sky130_fd_sc_hd__mux2_1 _10129_ (.A0(_05460_),
    .A1(\data_array.data0[11][20] ),
    .S(_03128_),
    .X(_01877_));
 sky130_fd_sc_hd__mux2_1 _10130_ (.A0(_05462_),
    .A1(\data_array.data0[11][21] ),
    .S(_03128_),
    .X(_01878_));
 sky130_fd_sc_hd__mux2_1 _10131_ (.A0(_05464_),
    .A1(\data_array.data0[11][22] ),
    .S(_03128_),
    .X(_01879_));
 sky130_fd_sc_hd__mux2_1 _10132_ (.A0(_05466_),
    .A1(\data_array.data0[11][23] ),
    .S(_03128_),
    .X(_01880_));
 sky130_fd_sc_hd__mux2_1 _10133_ (.A0(_05468_),
    .A1(\data_array.data0[11][24] ),
    .S(_03128_),
    .X(_01881_));
 sky130_fd_sc_hd__mux2_1 _10134_ (.A0(_05470_),
    .A1(\data_array.data0[11][25] ),
    .S(_03128_),
    .X(_01882_));
 sky130_fd_sc_hd__mux2_1 _10135_ (.A0(_05472_),
    .A1(\data_array.data0[11][26] ),
    .S(_03128_),
    .X(_01883_));
 sky130_fd_sc_hd__mux2_1 _10136_ (.A0(_05474_),
    .A1(\data_array.data0[11][27] ),
    .S(_03128_),
    .X(_01884_));
 sky130_fd_sc_hd__mux2_1 _10137_ (.A0(_05476_),
    .A1(\data_array.data0[11][28] ),
    .S(_03128_),
    .X(_01885_));
 sky130_fd_sc_hd__mux2_1 _10138_ (.A0(_05478_),
    .A1(\data_array.data0[11][29] ),
    .S(_03128_),
    .X(_01886_));
 sky130_fd_sc_hd__mux2_1 _10139_ (.A0(_05480_),
    .A1(\data_array.data0[11][30] ),
    .S(_03128_),
    .X(_01887_));
 sky130_fd_sc_hd__mux2_1 _10140_ (.A0(_05482_),
    .A1(\data_array.data0[11][31] ),
    .S(_03128_),
    .X(_01888_));
 sky130_fd_sc_hd__mux2_1 _10141_ (.A0(_05484_),
    .A1(\data_array.data0[11][32] ),
    .S(_03128_),
    .X(_01889_));
 sky130_fd_sc_hd__mux2_1 _10142_ (.A0(_05486_),
    .A1(\data_array.data0[11][33] ),
    .S(_03128_),
    .X(_01890_));
 sky130_fd_sc_hd__mux2_1 _10143_ (.A0(_05488_),
    .A1(\data_array.data0[11][34] ),
    .S(_03128_),
    .X(_01891_));
 sky130_fd_sc_hd__mux2_1 _10144_ (.A0(_05490_),
    .A1(\data_array.data0[11][35] ),
    .S(_03128_),
    .X(_01892_));
 sky130_fd_sc_hd__mux2_1 _10145_ (.A0(_05492_),
    .A1(\data_array.data0[11][36] ),
    .S(_03128_),
    .X(_01893_));
 sky130_fd_sc_hd__mux2_1 _10146_ (.A0(_05494_),
    .A1(\data_array.data0[11][37] ),
    .S(_03128_),
    .X(_01894_));
 sky130_fd_sc_hd__mux2_1 _10147_ (.A0(_05496_),
    .A1(\data_array.data0[11][38] ),
    .S(_03128_),
    .X(_01895_));
 sky130_fd_sc_hd__mux2_1 _10148_ (.A0(_05498_),
    .A1(\data_array.data0[11][39] ),
    .S(_03128_),
    .X(_01896_));
 sky130_fd_sc_hd__mux2_1 _10149_ (.A0(_05500_),
    .A1(\data_array.data0[11][40] ),
    .S(_03128_),
    .X(_01897_));
 sky130_fd_sc_hd__mux2_1 _10150_ (.A0(_05502_),
    .A1(\data_array.data0[11][41] ),
    .S(_03128_),
    .X(_01898_));
 sky130_fd_sc_hd__mux2_1 _10151_ (.A0(_05504_),
    .A1(\data_array.data0[11][42] ),
    .S(_03128_),
    .X(_01899_));
 sky130_fd_sc_hd__mux2_1 _10152_ (.A0(_05506_),
    .A1(\data_array.data0[11][43] ),
    .S(_03128_),
    .X(_01900_));
 sky130_fd_sc_hd__mux2_1 _10153_ (.A0(_05508_),
    .A1(\data_array.data0[11][44] ),
    .S(_03128_),
    .X(_01901_));
 sky130_fd_sc_hd__mux2_1 _10154_ (.A0(_05510_),
    .A1(\data_array.data0[11][45] ),
    .S(_03128_),
    .X(_01902_));
 sky130_fd_sc_hd__mux2_1 _10155_ (.A0(_05512_),
    .A1(\data_array.data0[11][46] ),
    .S(_03128_),
    .X(_01903_));
 sky130_fd_sc_hd__mux2_1 _10156_ (.A0(_05514_),
    .A1(\data_array.data0[11][47] ),
    .S(_03128_),
    .X(_01904_));
 sky130_fd_sc_hd__mux2_1 _10157_ (.A0(_05516_),
    .A1(\data_array.data0[11][48] ),
    .S(_03128_),
    .X(_01905_));
 sky130_fd_sc_hd__mux2_1 _10158_ (.A0(_05518_),
    .A1(\data_array.data0[11][49] ),
    .S(_03128_),
    .X(_01906_));
 sky130_fd_sc_hd__mux2_1 _10159_ (.A0(_05520_),
    .A1(\data_array.data0[11][50] ),
    .S(_03128_),
    .X(_01907_));
 sky130_fd_sc_hd__mux2_1 _10160_ (.A0(_05522_),
    .A1(\data_array.data0[11][51] ),
    .S(_03128_),
    .X(_01908_));
 sky130_fd_sc_hd__mux2_1 _10161_ (.A0(_05524_),
    .A1(\data_array.data0[11][52] ),
    .S(_03128_),
    .X(_01909_));
 sky130_fd_sc_hd__mux2_1 _10162_ (.A0(_05526_),
    .A1(\data_array.data0[11][53] ),
    .S(_03128_),
    .X(_01910_));
 sky130_fd_sc_hd__mux2_1 _10163_ (.A0(_05528_),
    .A1(\data_array.data0[11][54] ),
    .S(_03128_),
    .X(_01911_));
 sky130_fd_sc_hd__mux2_1 _10164_ (.A0(_05530_),
    .A1(\data_array.data0[11][55] ),
    .S(_03128_),
    .X(_01912_));
 sky130_fd_sc_hd__mux2_1 _10165_ (.A0(_05532_),
    .A1(\data_array.data0[11][56] ),
    .S(_03128_),
    .X(_01913_));
 sky130_fd_sc_hd__mux2_1 _10166_ (.A0(_05534_),
    .A1(\data_array.data0[11][57] ),
    .S(_03128_),
    .X(_01914_));
 sky130_fd_sc_hd__mux2_1 _10167_ (.A0(_05536_),
    .A1(\data_array.data0[11][58] ),
    .S(_03128_),
    .X(_01915_));
 sky130_fd_sc_hd__mux2_1 _10168_ (.A0(_05538_),
    .A1(\data_array.data0[11][59] ),
    .S(_03128_),
    .X(_01916_));
 sky130_fd_sc_hd__mux2_1 _10169_ (.A0(_05540_),
    .A1(\data_array.data0[11][60] ),
    .S(_03128_),
    .X(_01917_));
 sky130_fd_sc_hd__mux2_1 _10170_ (.A0(_05542_),
    .A1(\data_array.data0[11][61] ),
    .S(_03128_),
    .X(_01918_));
 sky130_fd_sc_hd__mux2_1 _10171_ (.A0(_05544_),
    .A1(\data_array.data0[11][62] ),
    .S(_03128_),
    .X(_01919_));
 sky130_fd_sc_hd__mux2_1 _10172_ (.A0(_05546_),
    .A1(\data_array.data0[11][63] ),
    .S(_03128_),
    .X(_01920_));
 sky130_fd_sc_hd__nand2_2 _10173_ (.A(_05415_),
    .B(_05547_),
    .Y(_03129_));
 sky130_fd_sc_hd__mux2_1 _10174_ (.A0(_05420_),
    .A1(\data_array.data0[10][0] ),
    .S(_03129_),
    .X(_01921_));
 sky130_fd_sc_hd__mux2_1 _10175_ (.A0(_05422_),
    .A1(\data_array.data0[10][1] ),
    .S(_03129_),
    .X(_01922_));
 sky130_fd_sc_hd__mux2_1 _10176_ (.A0(_05424_),
    .A1(\data_array.data0[10][2] ),
    .S(_03129_),
    .X(_01923_));
 sky130_fd_sc_hd__mux2_1 _10177_ (.A0(_05426_),
    .A1(\data_array.data0[10][3] ),
    .S(_03129_),
    .X(_01924_));
 sky130_fd_sc_hd__mux2_1 _10178_ (.A0(_05428_),
    .A1(\data_array.data0[10][4] ),
    .S(_03129_),
    .X(_01925_));
 sky130_fd_sc_hd__mux2_1 _10179_ (.A0(_05430_),
    .A1(\data_array.data0[10][5] ),
    .S(_03129_),
    .X(_01926_));
 sky130_fd_sc_hd__mux2_1 _10180_ (.A0(_05432_),
    .A1(\data_array.data0[10][6] ),
    .S(_03129_),
    .X(_01927_));
 sky130_fd_sc_hd__mux2_1 _10181_ (.A0(_05434_),
    .A1(\data_array.data0[10][7] ),
    .S(_03129_),
    .X(_01928_));
 sky130_fd_sc_hd__mux2_1 _10182_ (.A0(_05436_),
    .A1(\data_array.data0[10][8] ),
    .S(_03129_),
    .X(_01929_));
 sky130_fd_sc_hd__mux2_1 _10183_ (.A0(_05438_),
    .A1(\data_array.data0[10][9] ),
    .S(_03129_),
    .X(_01930_));
 sky130_fd_sc_hd__mux2_1 _10184_ (.A0(_05440_),
    .A1(\data_array.data0[10][10] ),
    .S(_03129_),
    .X(_01931_));
 sky130_fd_sc_hd__mux2_1 _10185_ (.A0(_05442_),
    .A1(\data_array.data0[10][11] ),
    .S(_03129_),
    .X(_01932_));
 sky130_fd_sc_hd__mux2_1 _10186_ (.A0(_05444_),
    .A1(\data_array.data0[10][12] ),
    .S(_03129_),
    .X(_01933_));
 sky130_fd_sc_hd__mux2_1 _10187_ (.A0(_05446_),
    .A1(\data_array.data0[10][13] ),
    .S(_03129_),
    .X(_01934_));
 sky130_fd_sc_hd__mux2_1 _10188_ (.A0(_05448_),
    .A1(\data_array.data0[10][14] ),
    .S(_03129_),
    .X(_01935_));
 sky130_fd_sc_hd__mux2_1 _10189_ (.A0(_05450_),
    .A1(\data_array.data0[10][15] ),
    .S(_03129_),
    .X(_01936_));
 sky130_fd_sc_hd__mux2_1 _10190_ (.A0(_05452_),
    .A1(\data_array.data0[10][16] ),
    .S(_03129_),
    .X(_01937_));
 sky130_fd_sc_hd__mux2_1 _10191_ (.A0(_05454_),
    .A1(\data_array.data0[10][17] ),
    .S(_03129_),
    .X(_01938_));
 sky130_fd_sc_hd__mux2_1 _10192_ (.A0(_05456_),
    .A1(\data_array.data0[10][18] ),
    .S(_03129_),
    .X(_01939_));
 sky130_fd_sc_hd__mux2_1 _10193_ (.A0(_05458_),
    .A1(\data_array.data0[10][19] ),
    .S(_03129_),
    .X(_01940_));
 sky130_fd_sc_hd__mux2_1 _10194_ (.A0(_05460_),
    .A1(\data_array.data0[10][20] ),
    .S(_03129_),
    .X(_01941_));
 sky130_fd_sc_hd__mux2_1 _10195_ (.A0(_05462_),
    .A1(\data_array.data0[10][21] ),
    .S(_03129_),
    .X(_01942_));
 sky130_fd_sc_hd__mux2_1 _10196_ (.A0(_05464_),
    .A1(\data_array.data0[10][22] ),
    .S(_03129_),
    .X(_01943_));
 sky130_fd_sc_hd__mux2_1 _10197_ (.A0(_05466_),
    .A1(\data_array.data0[10][23] ),
    .S(_03129_),
    .X(_01944_));
 sky130_fd_sc_hd__mux2_1 _10198_ (.A0(_05468_),
    .A1(\data_array.data0[10][24] ),
    .S(_03129_),
    .X(_01945_));
 sky130_fd_sc_hd__mux2_1 _10199_ (.A0(_05470_),
    .A1(\data_array.data0[10][25] ),
    .S(_03129_),
    .X(_01946_));
 sky130_fd_sc_hd__mux2_1 _10200_ (.A0(_05472_),
    .A1(\data_array.data0[10][26] ),
    .S(_03129_),
    .X(_01947_));
 sky130_fd_sc_hd__mux2_1 _10201_ (.A0(_05474_),
    .A1(\data_array.data0[10][27] ),
    .S(_03129_),
    .X(_01948_));
 sky130_fd_sc_hd__mux2_1 _10202_ (.A0(_05476_),
    .A1(\data_array.data0[10][28] ),
    .S(_03129_),
    .X(_01949_));
 sky130_fd_sc_hd__mux2_1 _10203_ (.A0(_05478_),
    .A1(\data_array.data0[10][29] ),
    .S(_03129_),
    .X(_01950_));
 sky130_fd_sc_hd__mux2_1 _10204_ (.A0(_05480_),
    .A1(\data_array.data0[10][30] ),
    .S(_03129_),
    .X(_01951_));
 sky130_fd_sc_hd__mux2_1 _10205_ (.A0(_05482_),
    .A1(\data_array.data0[10][31] ),
    .S(_03129_),
    .X(_01952_));
 sky130_fd_sc_hd__mux2_1 _10206_ (.A0(_05484_),
    .A1(\data_array.data0[10][32] ),
    .S(_03129_),
    .X(_01953_));
 sky130_fd_sc_hd__mux2_1 _10207_ (.A0(_05486_),
    .A1(\data_array.data0[10][33] ),
    .S(_03129_),
    .X(_01954_));
 sky130_fd_sc_hd__mux2_1 _10208_ (.A0(_05488_),
    .A1(\data_array.data0[10][34] ),
    .S(_03129_),
    .X(_01955_));
 sky130_fd_sc_hd__mux2_1 _10209_ (.A0(_05490_),
    .A1(\data_array.data0[10][35] ),
    .S(_03129_),
    .X(_01956_));
 sky130_fd_sc_hd__mux2_1 _10210_ (.A0(_05492_),
    .A1(\data_array.data0[10][36] ),
    .S(_03129_),
    .X(_01957_));
 sky130_fd_sc_hd__mux2_1 _10211_ (.A0(_05494_),
    .A1(\data_array.data0[10][37] ),
    .S(_03129_),
    .X(_01958_));
 sky130_fd_sc_hd__mux2_1 _10212_ (.A0(_05496_),
    .A1(\data_array.data0[10][38] ),
    .S(_03129_),
    .X(_01959_));
 sky130_fd_sc_hd__mux2_1 _10213_ (.A0(_05498_),
    .A1(\data_array.data0[10][39] ),
    .S(_03129_),
    .X(_01960_));
 sky130_fd_sc_hd__mux2_1 _10214_ (.A0(_05500_),
    .A1(\data_array.data0[10][40] ),
    .S(_03129_),
    .X(_01961_));
 sky130_fd_sc_hd__mux2_1 _10215_ (.A0(_05502_),
    .A1(\data_array.data0[10][41] ),
    .S(_03129_),
    .X(_01962_));
 sky130_fd_sc_hd__mux2_1 _10216_ (.A0(_05504_),
    .A1(\data_array.data0[10][42] ),
    .S(_03129_),
    .X(_01963_));
 sky130_fd_sc_hd__mux2_1 _10217_ (.A0(_05506_),
    .A1(\data_array.data0[10][43] ),
    .S(_03129_),
    .X(_01964_));
 sky130_fd_sc_hd__mux2_1 _10218_ (.A0(_05508_),
    .A1(\data_array.data0[10][44] ),
    .S(_03129_),
    .X(_01965_));
 sky130_fd_sc_hd__mux2_1 _10219_ (.A0(_05510_),
    .A1(\data_array.data0[10][45] ),
    .S(_03129_),
    .X(_01966_));
 sky130_fd_sc_hd__mux2_1 _10220_ (.A0(_05512_),
    .A1(\data_array.data0[10][46] ),
    .S(_03129_),
    .X(_01967_));
 sky130_fd_sc_hd__mux2_1 _10221_ (.A0(_05514_),
    .A1(\data_array.data0[10][47] ),
    .S(_03129_),
    .X(_01968_));
 sky130_fd_sc_hd__mux2_1 _10222_ (.A0(_05516_),
    .A1(\data_array.data0[10][48] ),
    .S(_03129_),
    .X(_01969_));
 sky130_fd_sc_hd__mux2_1 _10223_ (.A0(_05518_),
    .A1(\data_array.data0[10][49] ),
    .S(_03129_),
    .X(_01970_));
 sky130_fd_sc_hd__mux2_1 _10224_ (.A0(_05520_),
    .A1(\data_array.data0[10][50] ),
    .S(_03129_),
    .X(_01971_));
 sky130_fd_sc_hd__mux2_1 _10225_ (.A0(_05522_),
    .A1(\data_array.data0[10][51] ),
    .S(_03129_),
    .X(_01972_));
 sky130_fd_sc_hd__mux2_1 _10226_ (.A0(_05524_),
    .A1(\data_array.data0[10][52] ),
    .S(_03129_),
    .X(_01973_));
 sky130_fd_sc_hd__mux2_1 _10227_ (.A0(_05526_),
    .A1(\data_array.data0[10][53] ),
    .S(_03129_),
    .X(_01974_));
 sky130_fd_sc_hd__mux2_1 _10228_ (.A0(_05528_),
    .A1(\data_array.data0[10][54] ),
    .S(_03129_),
    .X(_01975_));
 sky130_fd_sc_hd__mux2_1 _10229_ (.A0(_05530_),
    .A1(\data_array.data0[10][55] ),
    .S(_03129_),
    .X(_01976_));
 sky130_fd_sc_hd__mux2_1 _10230_ (.A0(_05532_),
    .A1(\data_array.data0[10][56] ),
    .S(_03129_),
    .X(_01977_));
 sky130_fd_sc_hd__mux2_1 _10231_ (.A0(_05534_),
    .A1(\data_array.data0[10][57] ),
    .S(_03129_),
    .X(_01978_));
 sky130_fd_sc_hd__mux2_1 _10232_ (.A0(_05536_),
    .A1(\data_array.data0[10][58] ),
    .S(_03129_),
    .X(_01979_));
 sky130_fd_sc_hd__mux2_1 _10233_ (.A0(_05538_),
    .A1(\data_array.data0[10][59] ),
    .S(_03129_),
    .X(_01980_));
 sky130_fd_sc_hd__mux2_1 _10234_ (.A0(_05540_),
    .A1(\data_array.data0[10][60] ),
    .S(_03129_),
    .X(_01981_));
 sky130_fd_sc_hd__mux2_1 _10235_ (.A0(_05542_),
    .A1(\data_array.data0[10][61] ),
    .S(_03129_),
    .X(_01982_));
 sky130_fd_sc_hd__mux2_1 _10236_ (.A0(_05544_),
    .A1(\data_array.data0[10][62] ),
    .S(_03129_),
    .X(_01983_));
 sky130_fd_sc_hd__mux2_1 _10237_ (.A0(_05546_),
    .A1(\data_array.data0[10][63] ),
    .S(_03129_),
    .X(_01984_));
 sky130_fd_sc_hd__mux2_1 _10238_ (.A0(_05365_),
    .A1(\tag_array.tag0[2][0] ),
    .S(_05586_),
    .X(_01985_));
 sky130_fd_sc_hd__mux2_1 _10239_ (.A0(_05367_),
    .A1(\tag_array.tag0[2][1] ),
    .S(_05586_),
    .X(_01986_));
 sky130_fd_sc_hd__mux2_1 _10240_ (.A0(_05369_),
    .A1(\tag_array.tag0[2][2] ),
    .S(_05586_),
    .X(_01987_));
 sky130_fd_sc_hd__mux2_1 _10241_ (.A0(_05371_),
    .A1(\tag_array.tag0[2][3] ),
    .S(_05586_),
    .X(_01988_));
 sky130_fd_sc_hd__mux2_1 _10242_ (.A0(_05373_),
    .A1(\tag_array.tag0[2][4] ),
    .S(_05586_),
    .X(_01989_));
 sky130_fd_sc_hd__mux2_1 _10243_ (.A0(_05375_),
    .A1(\tag_array.tag0[2][5] ),
    .S(_05586_),
    .X(_01990_));
 sky130_fd_sc_hd__mux2_1 _10244_ (.A0(_05377_),
    .A1(\tag_array.tag0[2][6] ),
    .S(_05586_),
    .X(_01991_));
 sky130_fd_sc_hd__mux2_1 _10245_ (.A0(_05379_),
    .A1(\tag_array.tag0[2][7] ),
    .S(_05586_),
    .X(_01992_));
 sky130_fd_sc_hd__mux2_1 _10246_ (.A0(_05381_),
    .A1(\tag_array.tag0[2][8] ),
    .S(_05586_),
    .X(_01993_));
 sky130_fd_sc_hd__mux2_1 _10247_ (.A0(_05383_),
    .A1(\tag_array.tag0[2][9] ),
    .S(_05586_),
    .X(_01994_));
 sky130_fd_sc_hd__mux2_1 _10248_ (.A0(_05385_),
    .A1(\tag_array.tag0[2][10] ),
    .S(_05586_),
    .X(_01995_));
 sky130_fd_sc_hd__mux2_1 _10249_ (.A0(_05387_),
    .A1(\tag_array.tag0[2][11] ),
    .S(_05586_),
    .X(_01996_));
 sky130_fd_sc_hd__mux2_1 _10250_ (.A0(_05389_),
    .A1(\tag_array.tag0[2][12] ),
    .S(_05586_),
    .X(_01997_));
 sky130_fd_sc_hd__mux2_1 _10251_ (.A0(_05391_),
    .A1(\tag_array.tag0[2][13] ),
    .S(_05586_),
    .X(_01998_));
 sky130_fd_sc_hd__mux2_1 _10252_ (.A0(_05393_),
    .A1(\tag_array.tag0[2][14] ),
    .S(_05586_),
    .X(_01999_));
 sky130_fd_sc_hd__mux2_1 _10253_ (.A0(_05395_),
    .A1(\tag_array.tag0[2][15] ),
    .S(_05586_),
    .X(_02000_));
 sky130_fd_sc_hd__mux2_1 _10254_ (.A0(_05397_),
    .A1(\tag_array.tag0[2][16] ),
    .S(_05586_),
    .X(_02001_));
 sky130_fd_sc_hd__mux2_1 _10255_ (.A0(_05399_),
    .A1(\tag_array.tag0[2][17] ),
    .S(_05586_),
    .X(_02002_));
 sky130_fd_sc_hd__mux2_1 _10256_ (.A0(_05401_),
    .A1(\tag_array.tag0[2][18] ),
    .S(_05586_),
    .X(_02003_));
 sky130_fd_sc_hd__mux2_1 _10257_ (.A0(_05403_),
    .A1(\tag_array.tag0[2][19] ),
    .S(_05586_),
    .X(_02004_));
 sky130_fd_sc_hd__mux2_1 _10258_ (.A0(_05405_),
    .A1(\tag_array.tag0[2][20] ),
    .S(_05586_),
    .X(_02005_));
 sky130_fd_sc_hd__mux2_1 _10259_ (.A0(_05407_),
    .A1(\tag_array.tag0[2][21] ),
    .S(_05586_),
    .X(_02006_));
 sky130_fd_sc_hd__mux2_1 _10260_ (.A0(_05409_),
    .A1(\tag_array.tag0[2][22] ),
    .S(_05586_),
    .X(_02007_));
 sky130_fd_sc_hd__mux2_1 _10261_ (.A0(_05411_),
    .A1(\tag_array.tag0[2][23] ),
    .S(_05586_),
    .X(_02008_));
 sky130_fd_sc_hd__mux2_1 _10262_ (.A0(_05413_),
    .A1(\tag_array.tag0[2][24] ),
    .S(_05586_),
    .X(_02009_));
 sky130_fd_sc_hd__mux2_1 _10263_ (.A0(\data_array.data1[8][0] ),
    .A1(_05420_),
    .S(_05557_),
    .X(_02010_));
 sky130_fd_sc_hd__mux2_1 _10264_ (.A0(\data_array.data1[8][1] ),
    .A1(_05422_),
    .S(_05557_),
    .X(_02011_));
 sky130_fd_sc_hd__mux2_1 _10265_ (.A0(\data_array.data1[8][2] ),
    .A1(_05424_),
    .S(_05557_),
    .X(_02012_));
 sky130_fd_sc_hd__mux2_1 _10266_ (.A0(\data_array.data1[8][3] ),
    .A1(_05426_),
    .S(_05557_),
    .X(_02013_));
 sky130_fd_sc_hd__mux2_1 _10267_ (.A0(\data_array.data1[8][4] ),
    .A1(_05428_),
    .S(_05557_),
    .X(_02014_));
 sky130_fd_sc_hd__mux2_1 _10268_ (.A0(\data_array.data1[8][5] ),
    .A1(_05430_),
    .S(_05557_),
    .X(_02015_));
 sky130_fd_sc_hd__mux2_1 _10269_ (.A0(\data_array.data1[8][6] ),
    .A1(_05432_),
    .S(_05557_),
    .X(_02016_));
 sky130_fd_sc_hd__mux2_1 _10270_ (.A0(\data_array.data1[8][7] ),
    .A1(_05434_),
    .S(_05557_),
    .X(_02017_));
 sky130_fd_sc_hd__mux2_1 _10271_ (.A0(\data_array.data1[8][8] ),
    .A1(_05436_),
    .S(_05557_),
    .X(_02018_));
 sky130_fd_sc_hd__mux2_1 _10272_ (.A0(\data_array.data1[8][9] ),
    .A1(_05438_),
    .S(_05557_),
    .X(_02019_));
 sky130_fd_sc_hd__mux2_1 _10273_ (.A0(\data_array.data1[8][10] ),
    .A1(_05440_),
    .S(_05557_),
    .X(_02020_));
 sky130_fd_sc_hd__mux2_1 _10274_ (.A0(\data_array.data1[8][11] ),
    .A1(_05442_),
    .S(_05557_),
    .X(_02021_));
 sky130_fd_sc_hd__mux2_1 _10275_ (.A0(\data_array.data1[8][12] ),
    .A1(_05444_),
    .S(_05557_),
    .X(_02022_));
 sky130_fd_sc_hd__mux2_1 _10276_ (.A0(\data_array.data1[8][13] ),
    .A1(_05446_),
    .S(_05557_),
    .X(_02023_));
 sky130_fd_sc_hd__mux2_1 _10277_ (.A0(\data_array.data1[8][14] ),
    .A1(_05448_),
    .S(_05557_),
    .X(_02024_));
 sky130_fd_sc_hd__mux2_1 _10278_ (.A0(\data_array.data1[8][15] ),
    .A1(_05450_),
    .S(_05557_),
    .X(_02025_));
 sky130_fd_sc_hd__mux2_1 _10279_ (.A0(\data_array.data1[8][16] ),
    .A1(_05452_),
    .S(_05557_),
    .X(_02026_));
 sky130_fd_sc_hd__mux2_1 _10280_ (.A0(\data_array.data1[8][17] ),
    .A1(_05454_),
    .S(_05557_),
    .X(_02027_));
 sky130_fd_sc_hd__mux2_1 _10281_ (.A0(\data_array.data1[8][18] ),
    .A1(_05456_),
    .S(_05557_),
    .X(_02028_));
 sky130_fd_sc_hd__mux2_1 _10282_ (.A0(\data_array.data1[8][19] ),
    .A1(_05458_),
    .S(_05557_),
    .X(_02029_));
 sky130_fd_sc_hd__mux2_1 _10283_ (.A0(\data_array.data1[8][20] ),
    .A1(_05460_),
    .S(_05557_),
    .X(_02030_));
 sky130_fd_sc_hd__mux2_1 _10284_ (.A0(\data_array.data1[8][21] ),
    .A1(_05462_),
    .S(_05557_),
    .X(_02031_));
 sky130_fd_sc_hd__mux2_1 _10285_ (.A0(\data_array.data1[8][22] ),
    .A1(_05464_),
    .S(_05557_),
    .X(_02032_));
 sky130_fd_sc_hd__mux2_1 _10286_ (.A0(\data_array.data1[8][23] ),
    .A1(_05466_),
    .S(_05557_),
    .X(_02033_));
 sky130_fd_sc_hd__mux2_1 _10287_ (.A0(\data_array.data1[8][24] ),
    .A1(_05468_),
    .S(_05557_),
    .X(_02034_));
 sky130_fd_sc_hd__mux2_1 _10288_ (.A0(\data_array.data1[8][25] ),
    .A1(_05470_),
    .S(_05557_),
    .X(_02035_));
 sky130_fd_sc_hd__mux2_1 _10289_ (.A0(\data_array.data1[8][26] ),
    .A1(_05472_),
    .S(_05557_),
    .X(_02036_));
 sky130_fd_sc_hd__mux2_1 _10290_ (.A0(\data_array.data1[8][27] ),
    .A1(_05474_),
    .S(_05557_),
    .X(_02037_));
 sky130_fd_sc_hd__mux2_1 _10291_ (.A0(\data_array.data1[8][28] ),
    .A1(_05476_),
    .S(_05557_),
    .X(_02038_));
 sky130_fd_sc_hd__mux2_1 _10292_ (.A0(\data_array.data1[8][29] ),
    .A1(_05478_),
    .S(_05557_),
    .X(_02039_));
 sky130_fd_sc_hd__mux2_1 _10293_ (.A0(\data_array.data1[8][30] ),
    .A1(_05480_),
    .S(_05557_),
    .X(_02040_));
 sky130_fd_sc_hd__mux2_1 _10294_ (.A0(\data_array.data1[8][31] ),
    .A1(_05482_),
    .S(_05557_),
    .X(_02041_));
 sky130_fd_sc_hd__mux2_1 _10295_ (.A0(\data_array.data1[8][32] ),
    .A1(_05484_),
    .S(_05557_),
    .X(_02042_));
 sky130_fd_sc_hd__mux2_1 _10296_ (.A0(\data_array.data1[8][33] ),
    .A1(_05486_),
    .S(_05557_),
    .X(_02043_));
 sky130_fd_sc_hd__mux2_1 _10297_ (.A0(\data_array.data1[8][34] ),
    .A1(_05488_),
    .S(_05557_),
    .X(_02044_));
 sky130_fd_sc_hd__mux2_1 _10298_ (.A0(\data_array.data1[8][35] ),
    .A1(_05490_),
    .S(_05557_),
    .X(_02045_));
 sky130_fd_sc_hd__mux2_1 _10299_ (.A0(\data_array.data1[8][36] ),
    .A1(_05492_),
    .S(_05557_),
    .X(_02046_));
 sky130_fd_sc_hd__mux2_1 _10300_ (.A0(\data_array.data1[8][37] ),
    .A1(_05494_),
    .S(_05557_),
    .X(_02047_));
 sky130_fd_sc_hd__mux2_1 _10301_ (.A0(\data_array.data1[8][38] ),
    .A1(_05496_),
    .S(_05557_),
    .X(_02048_));
 sky130_fd_sc_hd__mux2_1 _10302_ (.A0(\data_array.data1[8][39] ),
    .A1(_05498_),
    .S(_05557_),
    .X(_02049_));
 sky130_fd_sc_hd__mux2_1 _10303_ (.A0(\data_array.data1[8][40] ),
    .A1(_05500_),
    .S(_05557_),
    .X(_02050_));
 sky130_fd_sc_hd__mux2_1 _10304_ (.A0(\data_array.data1[8][41] ),
    .A1(_05502_),
    .S(_05557_),
    .X(_02051_));
 sky130_fd_sc_hd__mux2_1 _10305_ (.A0(\data_array.data1[8][42] ),
    .A1(_05504_),
    .S(_05557_),
    .X(_02052_));
 sky130_fd_sc_hd__mux2_1 _10306_ (.A0(\data_array.data1[8][43] ),
    .A1(_05506_),
    .S(_05557_),
    .X(_02053_));
 sky130_fd_sc_hd__mux2_1 _10307_ (.A0(\data_array.data1[8][44] ),
    .A1(_05508_),
    .S(_05557_),
    .X(_02054_));
 sky130_fd_sc_hd__mux2_1 _10308_ (.A0(\data_array.data1[8][45] ),
    .A1(_05510_),
    .S(_05557_),
    .X(_02055_));
 sky130_fd_sc_hd__mux2_1 _10309_ (.A0(\data_array.data1[8][46] ),
    .A1(_05512_),
    .S(_05557_),
    .X(_02056_));
 sky130_fd_sc_hd__mux2_1 _10310_ (.A0(\data_array.data1[8][47] ),
    .A1(_05514_),
    .S(_05557_),
    .X(_02057_));
 sky130_fd_sc_hd__mux2_1 _10311_ (.A0(\data_array.data1[8][48] ),
    .A1(_05516_),
    .S(_05557_),
    .X(_02058_));
 sky130_fd_sc_hd__mux2_1 _10312_ (.A0(\data_array.data1[8][49] ),
    .A1(_05518_),
    .S(_05557_),
    .X(_02059_));
 sky130_fd_sc_hd__mux2_1 _10313_ (.A0(\data_array.data1[8][50] ),
    .A1(_05520_),
    .S(_05557_),
    .X(_02060_));
 sky130_fd_sc_hd__mux2_1 _10314_ (.A0(\data_array.data1[8][51] ),
    .A1(_05522_),
    .S(_05557_),
    .X(_02061_));
 sky130_fd_sc_hd__mux2_1 _10315_ (.A0(\data_array.data1[8][52] ),
    .A1(_05524_),
    .S(_05557_),
    .X(_02062_));
 sky130_fd_sc_hd__mux2_1 _10316_ (.A0(\data_array.data1[8][53] ),
    .A1(_05526_),
    .S(_05557_),
    .X(_02063_));
 sky130_fd_sc_hd__mux2_1 _10317_ (.A0(\data_array.data1[8][54] ),
    .A1(_05528_),
    .S(_05557_),
    .X(_02064_));
 sky130_fd_sc_hd__mux2_1 _10318_ (.A0(\data_array.data1[8][55] ),
    .A1(_05530_),
    .S(_05557_),
    .X(_02065_));
 sky130_fd_sc_hd__mux2_1 _10319_ (.A0(\data_array.data1[8][56] ),
    .A1(_05532_),
    .S(_05557_),
    .X(_02066_));
 sky130_fd_sc_hd__mux2_1 _10320_ (.A0(\data_array.data1[8][57] ),
    .A1(_05534_),
    .S(_05557_),
    .X(_02067_));
 sky130_fd_sc_hd__mux2_1 _10321_ (.A0(\data_array.data1[8][58] ),
    .A1(_05536_),
    .S(_05557_),
    .X(_02068_));
 sky130_fd_sc_hd__mux2_1 _10322_ (.A0(\data_array.data1[8][59] ),
    .A1(_05538_),
    .S(_05557_),
    .X(_02069_));
 sky130_fd_sc_hd__mux2_1 _10323_ (.A0(\data_array.data1[8][60] ),
    .A1(_05540_),
    .S(_05557_),
    .X(_02070_));
 sky130_fd_sc_hd__mux2_1 _10324_ (.A0(\data_array.data1[8][61] ),
    .A1(_05542_),
    .S(_05557_),
    .X(_02071_));
 sky130_fd_sc_hd__mux2_1 _10325_ (.A0(\data_array.data1[8][62] ),
    .A1(_05544_),
    .S(_05557_),
    .X(_02072_));
 sky130_fd_sc_hd__mux2_1 _10326_ (.A0(\data_array.data1[8][63] ),
    .A1(_05546_),
    .S(_05557_),
    .X(_02073_));
 sky130_fd_sc_hd__mux2_1 _10327_ (.A0(_05365_),
    .A1(\tag_array.tag0[1][0] ),
    .S(_05589_),
    .X(_02074_));
 sky130_fd_sc_hd__mux2_1 _10328_ (.A0(_05367_),
    .A1(\tag_array.tag0[1][1] ),
    .S(_05589_),
    .X(_02075_));
 sky130_fd_sc_hd__mux2_1 _10329_ (.A0(_05369_),
    .A1(\tag_array.tag0[1][2] ),
    .S(_05589_),
    .X(_02076_));
 sky130_fd_sc_hd__mux2_1 _10330_ (.A0(_05371_),
    .A1(\tag_array.tag0[1][3] ),
    .S(_05589_),
    .X(_02077_));
 sky130_fd_sc_hd__mux2_1 _10331_ (.A0(_05373_),
    .A1(\tag_array.tag0[1][4] ),
    .S(_05589_),
    .X(_02078_));
 sky130_fd_sc_hd__mux2_1 _10332_ (.A0(_05375_),
    .A1(\tag_array.tag0[1][5] ),
    .S(_05589_),
    .X(_02079_));
 sky130_fd_sc_hd__mux2_1 _10333_ (.A0(_05377_),
    .A1(\tag_array.tag0[1][6] ),
    .S(_05589_),
    .X(_02080_));
 sky130_fd_sc_hd__mux2_1 _10334_ (.A0(_05379_),
    .A1(\tag_array.tag0[1][7] ),
    .S(_05589_),
    .X(_02081_));
 sky130_fd_sc_hd__mux2_1 _10335_ (.A0(_05381_),
    .A1(\tag_array.tag0[1][8] ),
    .S(_05589_),
    .X(_02082_));
 sky130_fd_sc_hd__mux2_1 _10336_ (.A0(_05383_),
    .A1(\tag_array.tag0[1][9] ),
    .S(_05589_),
    .X(_02083_));
 sky130_fd_sc_hd__mux2_1 _10337_ (.A0(_05385_),
    .A1(\tag_array.tag0[1][10] ),
    .S(_05589_),
    .X(_02084_));
 sky130_fd_sc_hd__mux2_1 _10338_ (.A0(_05387_),
    .A1(\tag_array.tag0[1][11] ),
    .S(_05589_),
    .X(_02085_));
 sky130_fd_sc_hd__mux2_1 _10339_ (.A0(_05389_),
    .A1(\tag_array.tag0[1][12] ),
    .S(_05589_),
    .X(_02086_));
 sky130_fd_sc_hd__mux2_1 _10340_ (.A0(_05391_),
    .A1(\tag_array.tag0[1][13] ),
    .S(_05589_),
    .X(_02087_));
 sky130_fd_sc_hd__mux2_1 _10341_ (.A0(_05393_),
    .A1(\tag_array.tag0[1][14] ),
    .S(_05589_),
    .X(_02088_));
 sky130_fd_sc_hd__mux2_1 _10342_ (.A0(_05395_),
    .A1(\tag_array.tag0[1][15] ),
    .S(_05589_),
    .X(_02089_));
 sky130_fd_sc_hd__mux2_1 _10343_ (.A0(_05397_),
    .A1(\tag_array.tag0[1][16] ),
    .S(_05589_),
    .X(_02090_));
 sky130_fd_sc_hd__mux2_1 _10344_ (.A0(_05399_),
    .A1(\tag_array.tag0[1][17] ),
    .S(_05589_),
    .X(_02091_));
 sky130_fd_sc_hd__mux2_1 _10345_ (.A0(_05401_),
    .A1(\tag_array.tag0[1][18] ),
    .S(_05589_),
    .X(_02092_));
 sky130_fd_sc_hd__mux2_1 _10346_ (.A0(_05403_),
    .A1(\tag_array.tag0[1][19] ),
    .S(_05589_),
    .X(_02093_));
 sky130_fd_sc_hd__mux2_1 _10347_ (.A0(_05405_),
    .A1(\tag_array.tag0[1][20] ),
    .S(_05589_),
    .X(_02094_));
 sky130_fd_sc_hd__mux2_1 _10348_ (.A0(_05407_),
    .A1(\tag_array.tag0[1][21] ),
    .S(_05589_),
    .X(_02095_));
 sky130_fd_sc_hd__mux2_1 _10349_ (.A0(_05409_),
    .A1(\tag_array.tag0[1][22] ),
    .S(_05589_),
    .X(_02096_));
 sky130_fd_sc_hd__mux2_1 _10350_ (.A0(_05411_),
    .A1(\tag_array.tag0[1][23] ),
    .S(_05589_),
    .X(_02097_));
 sky130_fd_sc_hd__mux2_1 _10351_ (.A0(_05413_),
    .A1(\tag_array.tag0[1][24] ),
    .S(_05589_),
    .X(_02098_));
 sky130_fd_sc_hd__mux2_1 _10352_ (.A0(_05365_),
    .A1(\tag_array.tag0[15][0] ),
    .S(_05597_),
    .X(_02099_));
 sky130_fd_sc_hd__mux2_1 _10353_ (.A0(_05367_),
    .A1(\tag_array.tag0[15][1] ),
    .S(_05597_),
    .X(_02100_));
 sky130_fd_sc_hd__mux2_1 _10354_ (.A0(_05369_),
    .A1(\tag_array.tag0[15][2] ),
    .S(_05597_),
    .X(_02101_));
 sky130_fd_sc_hd__mux2_1 _10355_ (.A0(_05371_),
    .A1(\tag_array.tag0[15][3] ),
    .S(_05597_),
    .X(_02102_));
 sky130_fd_sc_hd__mux2_1 _10356_ (.A0(_05373_),
    .A1(\tag_array.tag0[15][4] ),
    .S(_05597_),
    .X(_02103_));
 sky130_fd_sc_hd__mux2_1 _10357_ (.A0(_05375_),
    .A1(\tag_array.tag0[15][5] ),
    .S(_05597_),
    .X(_02104_));
 sky130_fd_sc_hd__mux2_1 _10358_ (.A0(_05377_),
    .A1(\tag_array.tag0[15][6] ),
    .S(_05597_),
    .X(_02105_));
 sky130_fd_sc_hd__mux2_1 _10359_ (.A0(_05379_),
    .A1(\tag_array.tag0[15][7] ),
    .S(_05597_),
    .X(_02106_));
 sky130_fd_sc_hd__mux2_1 _10360_ (.A0(_05381_),
    .A1(\tag_array.tag0[15][8] ),
    .S(_05597_),
    .X(_02107_));
 sky130_fd_sc_hd__mux2_1 _10361_ (.A0(_05383_),
    .A1(\tag_array.tag0[15][9] ),
    .S(_05597_),
    .X(_02108_));
 sky130_fd_sc_hd__mux2_1 _10362_ (.A0(_05385_),
    .A1(\tag_array.tag0[15][10] ),
    .S(_05597_),
    .X(_02109_));
 sky130_fd_sc_hd__mux2_1 _10363_ (.A0(_05387_),
    .A1(\tag_array.tag0[15][11] ),
    .S(_05597_),
    .X(_02110_));
 sky130_fd_sc_hd__mux2_1 _10364_ (.A0(_05389_),
    .A1(\tag_array.tag0[15][12] ),
    .S(_05597_),
    .X(_02111_));
 sky130_fd_sc_hd__mux2_1 _10365_ (.A0(_05391_),
    .A1(\tag_array.tag0[15][13] ),
    .S(_05597_),
    .X(_02112_));
 sky130_fd_sc_hd__mux2_1 _10366_ (.A0(_05393_),
    .A1(\tag_array.tag0[15][14] ),
    .S(_05597_),
    .X(_02113_));
 sky130_fd_sc_hd__mux2_1 _10367_ (.A0(_05395_),
    .A1(\tag_array.tag0[15][15] ),
    .S(_05597_),
    .X(_02114_));
 sky130_fd_sc_hd__mux2_1 _10368_ (.A0(_05397_),
    .A1(\tag_array.tag0[15][16] ),
    .S(_05597_),
    .X(_02115_));
 sky130_fd_sc_hd__mux2_1 _10369_ (.A0(_05399_),
    .A1(\tag_array.tag0[15][17] ),
    .S(_05597_),
    .X(_02116_));
 sky130_fd_sc_hd__mux2_1 _10370_ (.A0(_05401_),
    .A1(\tag_array.tag0[15][18] ),
    .S(_05597_),
    .X(_02117_));
 sky130_fd_sc_hd__mux2_1 _10371_ (.A0(_05403_),
    .A1(\tag_array.tag0[15][19] ),
    .S(_05597_),
    .X(_02118_));
 sky130_fd_sc_hd__mux2_1 _10372_ (.A0(_05405_),
    .A1(\tag_array.tag0[15][20] ),
    .S(_05597_),
    .X(_02119_));
 sky130_fd_sc_hd__mux2_1 _10373_ (.A0(_05407_),
    .A1(\tag_array.tag0[15][21] ),
    .S(_05597_),
    .X(_02120_));
 sky130_fd_sc_hd__mux2_1 _10374_ (.A0(_05409_),
    .A1(\tag_array.tag0[15][22] ),
    .S(_05597_),
    .X(_02121_));
 sky130_fd_sc_hd__mux2_1 _10375_ (.A0(_05411_),
    .A1(\tag_array.tag0[15][23] ),
    .S(_05597_),
    .X(_02122_));
 sky130_fd_sc_hd__mux2_1 _10376_ (.A0(_05413_),
    .A1(\tag_array.tag0[15][24] ),
    .S(_05597_),
    .X(_02123_));
 sky130_fd_sc_hd__and2b_2 _10377_ (.A_N(_05353_),
    .B(cpu_write),
    .X(_03130_));
 sky130_fd_sc_hd__mux2_1 _10378_ (.A0(_03130_),
    .A1(\tag_array.dirty1[9] ),
    .S(_05591_),
    .X(_02124_));
 sky130_fd_sc_hd__mux2_1 _10379_ (.A0(_03130_),
    .A1(\tag_array.dirty1[14] ),
    .S(_05592_),
    .X(_02125_));
 sky130_fd_sc_hd__mux2_1 _10380_ (.A0(_03130_),
    .A1(\tag_array.dirty1[13] ),
    .S(_05593_),
    .X(_02126_));
 sky130_fd_sc_hd__mux2_1 _10381_ (.A0(_03130_),
    .A1(\tag_array.dirty1[12] ),
    .S(_05594_),
    .X(_02127_));
 sky130_fd_sc_hd__mux2_1 _10382_ (.A0(_03130_),
    .A1(\tag_array.dirty1[11] ),
    .S(_05551_),
    .X(_02128_));
 sky130_fd_sc_hd__mux2_1 _10383_ (.A0(_03130_),
    .A1(\tag_array.dirty1[10] ),
    .S(_05548_),
    .X(_02129_));
 sky130_fd_sc_hd__mux2_1 _10384_ (.A0(\tag_array.dirty1[0] ),
    .A1(_03130_),
    .S(_05549_),
    .X(_02130_));
 sky130_fd_sc_hd__mux2_1 _10385_ (.A0(\tag_array.dirty1[8] ),
    .A1(_03130_),
    .S(_05557_),
    .X(_02131_));
 sky130_fd_sc_hd__mux2_1 _10386_ (.A0(\data_array.data1[0][0] ),
    .A1(_05420_),
    .S(_05549_),
    .X(_02132_));
 sky130_fd_sc_hd__mux2_1 _10387_ (.A0(\data_array.data1[0][1] ),
    .A1(_05422_),
    .S(_05549_),
    .X(_02133_));
 sky130_fd_sc_hd__mux2_1 _10388_ (.A0(\data_array.data1[0][2] ),
    .A1(_05424_),
    .S(_05549_),
    .X(_02134_));
 sky130_fd_sc_hd__mux2_1 _10389_ (.A0(\data_array.data1[0][3] ),
    .A1(_05426_),
    .S(_05549_),
    .X(_02135_));
 sky130_fd_sc_hd__mux2_1 _10390_ (.A0(\data_array.data1[0][4] ),
    .A1(_05428_),
    .S(_05549_),
    .X(_02136_));
 sky130_fd_sc_hd__mux2_1 _10391_ (.A0(\data_array.data1[0][5] ),
    .A1(_05430_),
    .S(_05549_),
    .X(_02137_));
 sky130_fd_sc_hd__mux2_1 _10392_ (.A0(\data_array.data1[0][6] ),
    .A1(_05432_),
    .S(_05549_),
    .X(_02138_));
 sky130_fd_sc_hd__mux2_1 _10393_ (.A0(\data_array.data1[0][7] ),
    .A1(_05434_),
    .S(_05549_),
    .X(_02139_));
 sky130_fd_sc_hd__mux2_1 _10394_ (.A0(\data_array.data1[0][8] ),
    .A1(_05436_),
    .S(_05549_),
    .X(_02140_));
 sky130_fd_sc_hd__mux2_1 _10395_ (.A0(\data_array.data1[0][9] ),
    .A1(_05438_),
    .S(_05549_),
    .X(_02141_));
 sky130_fd_sc_hd__mux2_1 _10396_ (.A0(\data_array.data1[0][10] ),
    .A1(_05440_),
    .S(_05549_),
    .X(_02142_));
 sky130_fd_sc_hd__mux2_1 _10397_ (.A0(\data_array.data1[0][11] ),
    .A1(_05442_),
    .S(_05549_),
    .X(_02143_));
 sky130_fd_sc_hd__mux2_1 _10398_ (.A0(\data_array.data1[0][12] ),
    .A1(_05444_),
    .S(_05549_),
    .X(_02144_));
 sky130_fd_sc_hd__mux2_1 _10399_ (.A0(\data_array.data1[0][13] ),
    .A1(_05446_),
    .S(_05549_),
    .X(_02145_));
 sky130_fd_sc_hd__mux2_1 _10400_ (.A0(\data_array.data1[0][14] ),
    .A1(_05448_),
    .S(_05549_),
    .X(_02146_));
 sky130_fd_sc_hd__mux2_1 _10401_ (.A0(\data_array.data1[0][15] ),
    .A1(_05450_),
    .S(_05549_),
    .X(_02147_));
 sky130_fd_sc_hd__mux2_1 _10402_ (.A0(\data_array.data1[0][16] ),
    .A1(_05452_),
    .S(_05549_),
    .X(_02148_));
 sky130_fd_sc_hd__mux2_1 _10403_ (.A0(\data_array.data1[0][17] ),
    .A1(_05454_),
    .S(_05549_),
    .X(_02149_));
 sky130_fd_sc_hd__mux2_1 _10404_ (.A0(\data_array.data1[0][18] ),
    .A1(_05456_),
    .S(_05549_),
    .X(_02150_));
 sky130_fd_sc_hd__mux2_1 _10405_ (.A0(\data_array.data1[0][19] ),
    .A1(_05458_),
    .S(_05549_),
    .X(_02151_));
 sky130_fd_sc_hd__mux2_1 _10406_ (.A0(\data_array.data1[0][20] ),
    .A1(_05460_),
    .S(_05549_),
    .X(_02152_));
 sky130_fd_sc_hd__mux2_1 _10407_ (.A0(\data_array.data1[0][21] ),
    .A1(_05462_),
    .S(_05549_),
    .X(_02153_));
 sky130_fd_sc_hd__mux2_1 _10408_ (.A0(\data_array.data1[0][22] ),
    .A1(_05464_),
    .S(_05549_),
    .X(_02154_));
 sky130_fd_sc_hd__mux2_1 _10409_ (.A0(\data_array.data1[0][23] ),
    .A1(_05466_),
    .S(_05549_),
    .X(_02155_));
 sky130_fd_sc_hd__mux2_1 _10410_ (.A0(\data_array.data1[0][24] ),
    .A1(_05468_),
    .S(_05549_),
    .X(_02156_));
 sky130_fd_sc_hd__mux2_1 _10411_ (.A0(\data_array.data1[0][25] ),
    .A1(_05470_),
    .S(_05549_),
    .X(_02157_));
 sky130_fd_sc_hd__mux2_1 _10412_ (.A0(\data_array.data1[0][26] ),
    .A1(_05472_),
    .S(_05549_),
    .X(_02158_));
 sky130_fd_sc_hd__mux2_1 _10413_ (.A0(\data_array.data1[0][27] ),
    .A1(_05474_),
    .S(_05549_),
    .X(_02159_));
 sky130_fd_sc_hd__mux2_1 _10414_ (.A0(\data_array.data1[0][28] ),
    .A1(_05476_),
    .S(_05549_),
    .X(_02160_));
 sky130_fd_sc_hd__mux2_1 _10415_ (.A0(\data_array.data1[0][29] ),
    .A1(_05478_),
    .S(_05549_),
    .X(_02161_));
 sky130_fd_sc_hd__mux2_1 _10416_ (.A0(\data_array.data1[0][30] ),
    .A1(_05480_),
    .S(_05549_),
    .X(_02162_));
 sky130_fd_sc_hd__mux2_1 _10417_ (.A0(\data_array.data1[0][31] ),
    .A1(_05482_),
    .S(_05549_),
    .X(_02163_));
 sky130_fd_sc_hd__mux2_1 _10418_ (.A0(\data_array.data1[0][32] ),
    .A1(_05484_),
    .S(_05549_),
    .X(_02164_));
 sky130_fd_sc_hd__mux2_1 _10419_ (.A0(\data_array.data1[0][33] ),
    .A1(_05486_),
    .S(_05549_),
    .X(_02165_));
 sky130_fd_sc_hd__mux2_1 _10420_ (.A0(\data_array.data1[0][34] ),
    .A1(_05488_),
    .S(_05549_),
    .X(_02166_));
 sky130_fd_sc_hd__mux2_1 _10421_ (.A0(\data_array.data1[0][35] ),
    .A1(_05490_),
    .S(_05549_),
    .X(_02167_));
 sky130_fd_sc_hd__mux2_1 _10422_ (.A0(\data_array.data1[0][36] ),
    .A1(_05492_),
    .S(_05549_),
    .X(_02168_));
 sky130_fd_sc_hd__mux2_1 _10423_ (.A0(\data_array.data1[0][37] ),
    .A1(_05494_),
    .S(_05549_),
    .X(_02169_));
 sky130_fd_sc_hd__mux2_1 _10424_ (.A0(\data_array.data1[0][38] ),
    .A1(_05496_),
    .S(_05549_),
    .X(_02170_));
 sky130_fd_sc_hd__mux2_1 _10425_ (.A0(\data_array.data1[0][39] ),
    .A1(_05498_),
    .S(_05549_),
    .X(_02171_));
 sky130_fd_sc_hd__mux2_1 _10426_ (.A0(\data_array.data1[0][40] ),
    .A1(_05500_),
    .S(_05549_),
    .X(_02172_));
 sky130_fd_sc_hd__mux2_1 _10427_ (.A0(\data_array.data1[0][41] ),
    .A1(_05502_),
    .S(_05549_),
    .X(_02173_));
 sky130_fd_sc_hd__mux2_1 _10428_ (.A0(\data_array.data1[0][42] ),
    .A1(_05504_),
    .S(_05549_),
    .X(_02174_));
 sky130_fd_sc_hd__mux2_1 _10429_ (.A0(\data_array.data1[0][43] ),
    .A1(_05506_),
    .S(_05549_),
    .X(_02175_));
 sky130_fd_sc_hd__mux2_1 _10430_ (.A0(\data_array.data1[0][44] ),
    .A1(_05508_),
    .S(_05549_),
    .X(_02176_));
 sky130_fd_sc_hd__mux2_1 _10431_ (.A0(\data_array.data1[0][45] ),
    .A1(_05510_),
    .S(_05549_),
    .X(_02177_));
 sky130_fd_sc_hd__mux2_1 _10432_ (.A0(\data_array.data1[0][46] ),
    .A1(_05512_),
    .S(_05549_),
    .X(_02178_));
 sky130_fd_sc_hd__mux2_1 _10433_ (.A0(\data_array.data1[0][47] ),
    .A1(_05514_),
    .S(_05549_),
    .X(_02179_));
 sky130_fd_sc_hd__mux2_1 _10434_ (.A0(\data_array.data1[0][48] ),
    .A1(_05516_),
    .S(_05549_),
    .X(_02180_));
 sky130_fd_sc_hd__mux2_1 _10435_ (.A0(\data_array.data1[0][49] ),
    .A1(_05518_),
    .S(_05549_),
    .X(_02181_));
 sky130_fd_sc_hd__mux2_1 _10436_ (.A0(\data_array.data1[0][50] ),
    .A1(_05520_),
    .S(_05549_),
    .X(_02182_));
 sky130_fd_sc_hd__mux2_1 _10437_ (.A0(\data_array.data1[0][51] ),
    .A1(_05522_),
    .S(_05549_),
    .X(_02183_));
 sky130_fd_sc_hd__mux2_1 _10438_ (.A0(\data_array.data1[0][52] ),
    .A1(_05524_),
    .S(_05549_),
    .X(_02184_));
 sky130_fd_sc_hd__mux2_1 _10439_ (.A0(\data_array.data1[0][53] ),
    .A1(_05526_),
    .S(_05549_),
    .X(_02185_));
 sky130_fd_sc_hd__mux2_1 _10440_ (.A0(\data_array.data1[0][54] ),
    .A1(_05528_),
    .S(_05549_),
    .X(_02186_));
 sky130_fd_sc_hd__mux2_1 _10441_ (.A0(\data_array.data1[0][55] ),
    .A1(_05530_),
    .S(_05549_),
    .X(_02187_));
 sky130_fd_sc_hd__mux2_1 _10442_ (.A0(\data_array.data1[0][56] ),
    .A1(_05532_),
    .S(_05549_),
    .X(_02188_));
 sky130_fd_sc_hd__mux2_1 _10443_ (.A0(\data_array.data1[0][57] ),
    .A1(_05534_),
    .S(_05549_),
    .X(_02189_));
 sky130_fd_sc_hd__mux2_1 _10444_ (.A0(\data_array.data1[0][58] ),
    .A1(_05536_),
    .S(_05549_),
    .X(_02190_));
 sky130_fd_sc_hd__mux2_1 _10445_ (.A0(\data_array.data1[0][59] ),
    .A1(_05538_),
    .S(_05549_),
    .X(_02191_));
 sky130_fd_sc_hd__mux2_1 _10446_ (.A0(\data_array.data1[0][60] ),
    .A1(_05540_),
    .S(_05549_),
    .X(_02192_));
 sky130_fd_sc_hd__mux2_1 _10447_ (.A0(\data_array.data1[0][61] ),
    .A1(_05542_),
    .S(_05549_),
    .X(_02193_));
 sky130_fd_sc_hd__mux2_1 _10448_ (.A0(\data_array.data1[0][62] ),
    .A1(_05544_),
    .S(_05549_),
    .X(_02194_));
 sky130_fd_sc_hd__mux2_1 _10449_ (.A0(\data_array.data1[0][63] ),
    .A1(_05546_),
    .S(_05549_),
    .X(_02195_));
 sky130_fd_sc_hd__mux2_1 _10450_ (.A0(_03130_),
    .A1(\tag_array.dirty1[7] ),
    .S(_05362_),
    .X(_02196_));
 sky130_fd_sc_hd__mux2_1 _10451_ (.A0(_03130_),
    .A1(\tag_array.dirty1[6] ),
    .S(_05598_),
    .X(_02197_));
 sky130_fd_sc_hd__mux2_1 _10452_ (.A0(_03130_),
    .A1(\tag_array.dirty1[5] ),
    .S(_05599_),
    .X(_02198_));
 sky130_fd_sc_hd__mux2_1 _10453_ (.A0(\tag_array.dirty1[4] ),
    .A1(_03130_),
    .S(_05600_),
    .X(_02199_));
 sky130_fd_sc_hd__mux2_1 _10454_ (.A0(_03130_),
    .A1(\tag_array.dirty1[3] ),
    .S(_05601_),
    .X(_02200_));
 sky130_fd_sc_hd__mux2_1 _10455_ (.A0(\tag_array.dirty1[2] ),
    .A1(_03130_),
    .S(_05602_),
    .X(_02201_));
 sky130_fd_sc_hd__mux2_1 _10456_ (.A0(\tag_array.dirty1[1] ),
    .A1(_03130_),
    .S(_05603_),
    .X(_02202_));
 sky130_fd_sc_hd__mux2_1 _10457_ (.A0(_03130_),
    .A1(\tag_array.dirty1[15] ),
    .S(_05604_),
    .X(_02203_));
 sky130_fd_sc_hd__nand2_2 _10458_ (.A(_05415_),
    .B(_05590_),
    .Y(_03131_));
 sky130_fd_sc_hd__mux2_1 _10459_ (.A0(_05420_),
    .A1(\data_array.data0[9][0] ),
    .S(_03131_),
    .X(_02204_));
 sky130_fd_sc_hd__mux2_1 _10460_ (.A0(_05422_),
    .A1(\data_array.data0[9][1] ),
    .S(_03131_),
    .X(_02205_));
 sky130_fd_sc_hd__mux2_1 _10461_ (.A0(_05424_),
    .A1(\data_array.data0[9][2] ),
    .S(_03131_),
    .X(_02206_));
 sky130_fd_sc_hd__mux2_1 _10462_ (.A0(_05426_),
    .A1(\data_array.data0[9][3] ),
    .S(_03131_),
    .X(_02207_));
 sky130_fd_sc_hd__mux2_1 _10463_ (.A0(_05428_),
    .A1(\data_array.data0[9][4] ),
    .S(_03131_),
    .X(_02208_));
 sky130_fd_sc_hd__mux2_1 _10464_ (.A0(_05430_),
    .A1(\data_array.data0[9][5] ),
    .S(_03131_),
    .X(_02209_));
 sky130_fd_sc_hd__mux2_1 _10465_ (.A0(_05432_),
    .A1(\data_array.data0[9][6] ),
    .S(_03131_),
    .X(_02210_));
 sky130_fd_sc_hd__mux2_1 _10466_ (.A0(_05434_),
    .A1(\data_array.data0[9][7] ),
    .S(_03131_),
    .X(_02211_));
 sky130_fd_sc_hd__mux2_1 _10467_ (.A0(_05436_),
    .A1(\data_array.data0[9][8] ),
    .S(_03131_),
    .X(_02212_));
 sky130_fd_sc_hd__mux2_1 _10468_ (.A0(_05438_),
    .A1(\data_array.data0[9][9] ),
    .S(_03131_),
    .X(_02213_));
 sky130_fd_sc_hd__mux2_1 _10469_ (.A0(_05440_),
    .A1(\data_array.data0[9][10] ),
    .S(_03131_),
    .X(_02214_));
 sky130_fd_sc_hd__mux2_1 _10470_ (.A0(_05442_),
    .A1(\data_array.data0[9][11] ),
    .S(_03131_),
    .X(_02215_));
 sky130_fd_sc_hd__mux2_1 _10471_ (.A0(_05444_),
    .A1(\data_array.data0[9][12] ),
    .S(_03131_),
    .X(_02216_));
 sky130_fd_sc_hd__mux2_1 _10472_ (.A0(_05446_),
    .A1(\data_array.data0[9][13] ),
    .S(_03131_),
    .X(_02217_));
 sky130_fd_sc_hd__mux2_1 _10473_ (.A0(_05448_),
    .A1(\data_array.data0[9][14] ),
    .S(_03131_),
    .X(_02218_));
 sky130_fd_sc_hd__mux2_1 _10474_ (.A0(_05450_),
    .A1(\data_array.data0[9][15] ),
    .S(_03131_),
    .X(_02219_));
 sky130_fd_sc_hd__mux2_1 _10475_ (.A0(_05452_),
    .A1(\data_array.data0[9][16] ),
    .S(_03131_),
    .X(_02220_));
 sky130_fd_sc_hd__mux2_1 _10476_ (.A0(_05454_),
    .A1(\data_array.data0[9][17] ),
    .S(_03131_),
    .X(_02221_));
 sky130_fd_sc_hd__mux2_1 _10477_ (.A0(_05456_),
    .A1(\data_array.data0[9][18] ),
    .S(_03131_),
    .X(_02222_));
 sky130_fd_sc_hd__mux2_1 _10478_ (.A0(_05458_),
    .A1(\data_array.data0[9][19] ),
    .S(_03131_),
    .X(_02223_));
 sky130_fd_sc_hd__mux2_1 _10479_ (.A0(_05460_),
    .A1(\data_array.data0[9][20] ),
    .S(_03131_),
    .X(_02224_));
 sky130_fd_sc_hd__mux2_1 _10480_ (.A0(_05462_),
    .A1(\data_array.data0[9][21] ),
    .S(_03131_),
    .X(_02225_));
 sky130_fd_sc_hd__mux2_1 _10481_ (.A0(_05464_),
    .A1(\data_array.data0[9][22] ),
    .S(_03131_),
    .X(_02226_));
 sky130_fd_sc_hd__mux2_1 _10482_ (.A0(_05466_),
    .A1(\data_array.data0[9][23] ),
    .S(_03131_),
    .X(_02227_));
 sky130_fd_sc_hd__mux2_1 _10483_ (.A0(_05468_),
    .A1(\data_array.data0[9][24] ),
    .S(_03131_),
    .X(_02228_));
 sky130_fd_sc_hd__mux2_1 _10484_ (.A0(_05470_),
    .A1(\data_array.data0[9][25] ),
    .S(_03131_),
    .X(_02229_));
 sky130_fd_sc_hd__mux2_1 _10485_ (.A0(_05472_),
    .A1(\data_array.data0[9][26] ),
    .S(_03131_),
    .X(_02230_));
 sky130_fd_sc_hd__mux2_1 _10486_ (.A0(_05474_),
    .A1(\data_array.data0[9][27] ),
    .S(_03131_),
    .X(_02231_));
 sky130_fd_sc_hd__mux2_1 _10487_ (.A0(_05476_),
    .A1(\data_array.data0[9][28] ),
    .S(_03131_),
    .X(_02232_));
 sky130_fd_sc_hd__mux2_1 _10488_ (.A0(_05478_),
    .A1(\data_array.data0[9][29] ),
    .S(_03131_),
    .X(_02233_));
 sky130_fd_sc_hd__mux2_1 _10489_ (.A0(_05480_),
    .A1(\data_array.data0[9][30] ),
    .S(_03131_),
    .X(_02234_));
 sky130_fd_sc_hd__mux2_1 _10490_ (.A0(_05482_),
    .A1(\data_array.data0[9][31] ),
    .S(_03131_),
    .X(_02235_));
 sky130_fd_sc_hd__mux2_1 _10491_ (.A0(_05484_),
    .A1(\data_array.data0[9][32] ),
    .S(_03131_),
    .X(_02236_));
 sky130_fd_sc_hd__mux2_1 _10492_ (.A0(_05486_),
    .A1(\data_array.data0[9][33] ),
    .S(_03131_),
    .X(_02237_));
 sky130_fd_sc_hd__mux2_1 _10493_ (.A0(_05488_),
    .A1(\data_array.data0[9][34] ),
    .S(_03131_),
    .X(_02238_));
 sky130_fd_sc_hd__mux2_1 _10494_ (.A0(_05490_),
    .A1(\data_array.data0[9][35] ),
    .S(_03131_),
    .X(_02239_));
 sky130_fd_sc_hd__mux2_1 _10495_ (.A0(_05492_),
    .A1(\data_array.data0[9][36] ),
    .S(_03131_),
    .X(_02240_));
 sky130_fd_sc_hd__mux2_1 _10496_ (.A0(_05494_),
    .A1(\data_array.data0[9][37] ),
    .S(_03131_),
    .X(_02241_));
 sky130_fd_sc_hd__mux2_1 _10497_ (.A0(_05496_),
    .A1(\data_array.data0[9][38] ),
    .S(_03131_),
    .X(_02242_));
 sky130_fd_sc_hd__mux2_1 _10498_ (.A0(_05498_),
    .A1(\data_array.data0[9][39] ),
    .S(_03131_),
    .X(_02243_));
 sky130_fd_sc_hd__mux2_1 _10499_ (.A0(_05500_),
    .A1(\data_array.data0[9][40] ),
    .S(_03131_),
    .X(_02244_));
 sky130_fd_sc_hd__mux2_1 _10500_ (.A0(_05502_),
    .A1(\data_array.data0[9][41] ),
    .S(_03131_),
    .X(_02245_));
 sky130_fd_sc_hd__mux2_1 _10501_ (.A0(_05504_),
    .A1(\data_array.data0[9][42] ),
    .S(_03131_),
    .X(_02246_));
 sky130_fd_sc_hd__mux2_1 _10502_ (.A0(_05506_),
    .A1(\data_array.data0[9][43] ),
    .S(_03131_),
    .X(_02247_));
 sky130_fd_sc_hd__mux2_1 _10503_ (.A0(_05508_),
    .A1(\data_array.data0[9][44] ),
    .S(_03131_),
    .X(_02248_));
 sky130_fd_sc_hd__mux2_1 _10504_ (.A0(_05510_),
    .A1(\data_array.data0[9][45] ),
    .S(_03131_),
    .X(_02249_));
 sky130_fd_sc_hd__mux2_1 _10505_ (.A0(_05512_),
    .A1(\data_array.data0[9][46] ),
    .S(_03131_),
    .X(_02250_));
 sky130_fd_sc_hd__mux2_1 _10506_ (.A0(_05514_),
    .A1(\data_array.data0[9][47] ),
    .S(_03131_),
    .X(_02251_));
 sky130_fd_sc_hd__mux2_1 _10507_ (.A0(_05516_),
    .A1(\data_array.data0[9][48] ),
    .S(_03131_),
    .X(_02252_));
 sky130_fd_sc_hd__mux2_1 _10508_ (.A0(_05518_),
    .A1(\data_array.data0[9][49] ),
    .S(_03131_),
    .X(_02253_));
 sky130_fd_sc_hd__mux2_1 _10509_ (.A0(_05520_),
    .A1(\data_array.data0[9][50] ),
    .S(_03131_),
    .X(_02254_));
 sky130_fd_sc_hd__mux2_1 _10510_ (.A0(_05522_),
    .A1(\data_array.data0[9][51] ),
    .S(_03131_),
    .X(_02255_));
 sky130_fd_sc_hd__mux2_1 _10511_ (.A0(_05524_),
    .A1(\data_array.data0[9][52] ),
    .S(_03131_),
    .X(_02256_));
 sky130_fd_sc_hd__mux2_1 _10512_ (.A0(_05526_),
    .A1(\data_array.data0[9][53] ),
    .S(_03131_),
    .X(_02257_));
 sky130_fd_sc_hd__mux2_1 _10513_ (.A0(_05528_),
    .A1(\data_array.data0[9][54] ),
    .S(_03131_),
    .X(_02258_));
 sky130_fd_sc_hd__mux2_1 _10514_ (.A0(_05530_),
    .A1(\data_array.data0[9][55] ),
    .S(_03131_),
    .X(_02259_));
 sky130_fd_sc_hd__mux2_1 _10515_ (.A0(_05532_),
    .A1(\data_array.data0[9][56] ),
    .S(_03131_),
    .X(_02260_));
 sky130_fd_sc_hd__mux2_1 _10516_ (.A0(_05534_),
    .A1(\data_array.data0[9][57] ),
    .S(_03131_),
    .X(_02261_));
 sky130_fd_sc_hd__mux2_1 _10517_ (.A0(_05536_),
    .A1(\data_array.data0[9][58] ),
    .S(_03131_),
    .X(_02262_));
 sky130_fd_sc_hd__mux2_1 _10518_ (.A0(_05538_),
    .A1(\data_array.data0[9][59] ),
    .S(_03131_),
    .X(_02263_));
 sky130_fd_sc_hd__mux2_1 _10519_ (.A0(_05540_),
    .A1(\data_array.data0[9][60] ),
    .S(_03131_),
    .X(_02264_));
 sky130_fd_sc_hd__mux2_1 _10520_ (.A0(_05542_),
    .A1(\data_array.data0[9][61] ),
    .S(_03131_),
    .X(_02265_));
 sky130_fd_sc_hd__mux2_1 _10521_ (.A0(_05544_),
    .A1(\data_array.data0[9][62] ),
    .S(_03131_),
    .X(_02266_));
 sky130_fd_sc_hd__mux2_1 _10522_ (.A0(_05546_),
    .A1(\data_array.data0[9][63] ),
    .S(_03131_),
    .X(_02267_));
 sky130_fd_sc_hd__mux2_1 _10523_ (.A0(cpu_write),
    .A1(\tag_array.dirty0[9] ),
    .S(_05606_),
    .X(_02268_));
 sky130_fd_sc_hd__mux2_1 _10524_ (.A0(_05420_),
    .A1(\data_array.data1[15][0] ),
    .S(_05604_),
    .X(_02269_));
 sky130_fd_sc_hd__mux2_1 _10525_ (.A0(_05422_),
    .A1(\data_array.data1[15][1] ),
    .S(_05604_),
    .X(_02270_));
 sky130_fd_sc_hd__mux2_1 _10526_ (.A0(_05424_),
    .A1(\data_array.data1[15][2] ),
    .S(_05604_),
    .X(_02271_));
 sky130_fd_sc_hd__mux2_1 _10527_ (.A0(_05426_),
    .A1(\data_array.data1[15][3] ),
    .S(_05604_),
    .X(_02272_));
 sky130_fd_sc_hd__mux2_1 _10528_ (.A0(_05428_),
    .A1(\data_array.data1[15][4] ),
    .S(_05604_),
    .X(_02273_));
 sky130_fd_sc_hd__mux2_1 _10529_ (.A0(_05430_),
    .A1(\data_array.data1[15][5] ),
    .S(_05604_),
    .X(_02274_));
 sky130_fd_sc_hd__mux2_1 _10530_ (.A0(_05432_),
    .A1(\data_array.data1[15][6] ),
    .S(_05604_),
    .X(_02275_));
 sky130_fd_sc_hd__mux2_1 _10531_ (.A0(_05434_),
    .A1(\data_array.data1[15][7] ),
    .S(_05604_),
    .X(_02276_));
 sky130_fd_sc_hd__mux2_1 _10532_ (.A0(_05436_),
    .A1(\data_array.data1[15][8] ),
    .S(_05604_),
    .X(_02277_));
 sky130_fd_sc_hd__mux2_1 _10533_ (.A0(_05438_),
    .A1(\data_array.data1[15][9] ),
    .S(_05604_),
    .X(_02278_));
 sky130_fd_sc_hd__mux2_1 _10534_ (.A0(_05440_),
    .A1(\data_array.data1[15][10] ),
    .S(_05604_),
    .X(_02279_));
 sky130_fd_sc_hd__mux2_1 _10535_ (.A0(_05442_),
    .A1(\data_array.data1[15][11] ),
    .S(_05604_),
    .X(_02280_));
 sky130_fd_sc_hd__mux2_1 _10536_ (.A0(_05444_),
    .A1(\data_array.data1[15][12] ),
    .S(_05604_),
    .X(_02281_));
 sky130_fd_sc_hd__mux2_1 _10537_ (.A0(_05446_),
    .A1(\data_array.data1[15][13] ),
    .S(_05604_),
    .X(_02282_));
 sky130_fd_sc_hd__mux2_1 _10538_ (.A0(_05448_),
    .A1(\data_array.data1[15][14] ),
    .S(_05604_),
    .X(_02283_));
 sky130_fd_sc_hd__mux2_1 _10539_ (.A0(_05450_),
    .A1(\data_array.data1[15][15] ),
    .S(_05604_),
    .X(_02284_));
 sky130_fd_sc_hd__mux2_1 _10540_ (.A0(_05452_),
    .A1(\data_array.data1[15][16] ),
    .S(_05604_),
    .X(_02285_));
 sky130_fd_sc_hd__mux2_1 _10541_ (.A0(_05454_),
    .A1(\data_array.data1[15][17] ),
    .S(_05604_),
    .X(_02286_));
 sky130_fd_sc_hd__mux2_1 _10542_ (.A0(_05456_),
    .A1(\data_array.data1[15][18] ),
    .S(_05604_),
    .X(_02287_));
 sky130_fd_sc_hd__mux2_1 _10543_ (.A0(_05458_),
    .A1(\data_array.data1[15][19] ),
    .S(_05604_),
    .X(_02288_));
 sky130_fd_sc_hd__mux2_1 _10544_ (.A0(_05460_),
    .A1(\data_array.data1[15][20] ),
    .S(_05604_),
    .X(_02289_));
 sky130_fd_sc_hd__mux2_1 _10545_ (.A0(_05462_),
    .A1(\data_array.data1[15][21] ),
    .S(_05604_),
    .X(_02290_));
 sky130_fd_sc_hd__mux2_1 _10546_ (.A0(_05464_),
    .A1(\data_array.data1[15][22] ),
    .S(_05604_),
    .X(_02291_));
 sky130_fd_sc_hd__mux2_1 _10547_ (.A0(_05466_),
    .A1(\data_array.data1[15][23] ),
    .S(_05604_),
    .X(_02292_));
 sky130_fd_sc_hd__mux2_1 _10548_ (.A0(_05468_),
    .A1(\data_array.data1[15][24] ),
    .S(_05604_),
    .X(_02293_));
 sky130_fd_sc_hd__mux2_1 _10549_ (.A0(_05470_),
    .A1(\data_array.data1[15][25] ),
    .S(_05604_),
    .X(_02294_));
 sky130_fd_sc_hd__mux2_1 _10550_ (.A0(_05472_),
    .A1(\data_array.data1[15][26] ),
    .S(_05604_),
    .X(_02295_));
 sky130_fd_sc_hd__mux2_1 _10551_ (.A0(_05474_),
    .A1(\data_array.data1[15][27] ),
    .S(_05604_),
    .X(_02296_));
 sky130_fd_sc_hd__mux2_1 _10552_ (.A0(_05476_),
    .A1(\data_array.data1[15][28] ),
    .S(_05604_),
    .X(_02297_));
 sky130_fd_sc_hd__mux2_1 _10553_ (.A0(_05478_),
    .A1(\data_array.data1[15][29] ),
    .S(_05604_),
    .X(_02298_));
 sky130_fd_sc_hd__mux2_1 _10554_ (.A0(_05480_),
    .A1(\data_array.data1[15][30] ),
    .S(_05604_),
    .X(_02299_));
 sky130_fd_sc_hd__mux2_1 _10555_ (.A0(_05482_),
    .A1(\data_array.data1[15][31] ),
    .S(_05604_),
    .X(_02300_));
 sky130_fd_sc_hd__mux2_1 _10556_ (.A0(_05484_),
    .A1(\data_array.data1[15][32] ),
    .S(_05604_),
    .X(_02301_));
 sky130_fd_sc_hd__mux2_1 _10557_ (.A0(_05486_),
    .A1(\data_array.data1[15][33] ),
    .S(_05604_),
    .X(_02302_));
 sky130_fd_sc_hd__mux2_1 _10558_ (.A0(_05488_),
    .A1(\data_array.data1[15][34] ),
    .S(_05604_),
    .X(_02303_));
 sky130_fd_sc_hd__mux2_1 _10559_ (.A0(_05490_),
    .A1(\data_array.data1[15][35] ),
    .S(_05604_),
    .X(_02304_));
 sky130_fd_sc_hd__mux2_1 _10560_ (.A0(_05492_),
    .A1(\data_array.data1[15][36] ),
    .S(_05604_),
    .X(_02305_));
 sky130_fd_sc_hd__mux2_1 _10561_ (.A0(_05494_),
    .A1(\data_array.data1[15][37] ),
    .S(_05604_),
    .X(_02306_));
 sky130_fd_sc_hd__mux2_1 _10562_ (.A0(_05496_),
    .A1(\data_array.data1[15][38] ),
    .S(_05604_),
    .X(_02307_));
 sky130_fd_sc_hd__mux2_1 _10563_ (.A0(_05498_),
    .A1(\data_array.data1[15][39] ),
    .S(_05604_),
    .X(_02308_));
 sky130_fd_sc_hd__mux2_1 _10564_ (.A0(_05500_),
    .A1(\data_array.data1[15][40] ),
    .S(_05604_),
    .X(_02309_));
 sky130_fd_sc_hd__mux2_1 _10565_ (.A0(_05502_),
    .A1(\data_array.data1[15][41] ),
    .S(_05604_),
    .X(_02310_));
 sky130_fd_sc_hd__mux2_1 _10566_ (.A0(_05504_),
    .A1(\data_array.data1[15][42] ),
    .S(_05604_),
    .X(_02311_));
 sky130_fd_sc_hd__mux2_1 _10567_ (.A0(_05506_),
    .A1(\data_array.data1[15][43] ),
    .S(_05604_),
    .X(_02312_));
 sky130_fd_sc_hd__mux2_1 _10568_ (.A0(_05508_),
    .A1(\data_array.data1[15][44] ),
    .S(_05604_),
    .X(_02313_));
 sky130_fd_sc_hd__mux2_1 _10569_ (.A0(_05510_),
    .A1(\data_array.data1[15][45] ),
    .S(_05604_),
    .X(_02314_));
 sky130_fd_sc_hd__mux2_1 _10570_ (.A0(_05512_),
    .A1(\data_array.data1[15][46] ),
    .S(_05604_),
    .X(_02315_));
 sky130_fd_sc_hd__mux2_1 _10571_ (.A0(_05514_),
    .A1(\data_array.data1[15][47] ),
    .S(_05604_),
    .X(_02316_));
 sky130_fd_sc_hd__mux2_1 _10572_ (.A0(_05516_),
    .A1(\data_array.data1[15][48] ),
    .S(_05604_),
    .X(_02317_));
 sky130_fd_sc_hd__mux2_1 _10573_ (.A0(_05518_),
    .A1(\data_array.data1[15][49] ),
    .S(_05604_),
    .X(_02318_));
 sky130_fd_sc_hd__mux2_1 _10574_ (.A0(_05520_),
    .A1(\data_array.data1[15][50] ),
    .S(_05604_),
    .X(_02319_));
 sky130_fd_sc_hd__mux2_1 _10575_ (.A0(_05522_),
    .A1(\data_array.data1[15][51] ),
    .S(_05604_),
    .X(_02320_));
 sky130_fd_sc_hd__mux2_1 _10576_ (.A0(_05524_),
    .A1(\data_array.data1[15][52] ),
    .S(_05604_),
    .X(_02321_));
 sky130_fd_sc_hd__mux2_1 _10577_ (.A0(_05526_),
    .A1(\data_array.data1[15][53] ),
    .S(_05604_),
    .X(_02322_));
 sky130_fd_sc_hd__mux2_1 _10578_ (.A0(_05528_),
    .A1(\data_array.data1[15][54] ),
    .S(_05604_),
    .X(_02323_));
 sky130_fd_sc_hd__mux2_1 _10579_ (.A0(_05530_),
    .A1(\data_array.data1[15][55] ),
    .S(_05604_),
    .X(_02324_));
 sky130_fd_sc_hd__mux2_1 _10580_ (.A0(_05532_),
    .A1(\data_array.data1[15][56] ),
    .S(_05604_),
    .X(_02325_));
 sky130_fd_sc_hd__mux2_1 _10581_ (.A0(_05534_),
    .A1(\data_array.data1[15][57] ),
    .S(_05604_),
    .X(_02326_));
 sky130_fd_sc_hd__mux2_1 _10582_ (.A0(_05536_),
    .A1(\data_array.data1[15][58] ),
    .S(_05604_),
    .X(_02327_));
 sky130_fd_sc_hd__mux2_1 _10583_ (.A0(_05538_),
    .A1(\data_array.data1[15][59] ),
    .S(_05604_),
    .X(_02328_));
 sky130_fd_sc_hd__mux2_1 _10584_ (.A0(_05540_),
    .A1(\data_array.data1[15][60] ),
    .S(_05604_),
    .X(_02329_));
 sky130_fd_sc_hd__mux2_1 _10585_ (.A0(_05542_),
    .A1(\data_array.data1[15][61] ),
    .S(_05604_),
    .X(_02330_));
 sky130_fd_sc_hd__mux2_1 _10586_ (.A0(_05544_),
    .A1(\data_array.data1[15][62] ),
    .S(_05604_),
    .X(_02331_));
 sky130_fd_sc_hd__mux2_1 _10587_ (.A0(_05546_),
    .A1(\data_array.data1[15][63] ),
    .S(_05604_),
    .X(_02332_));
 sky130_fd_sc_hd__mux2_1 _10588_ (.A0(\data_array.data1[1][0] ),
    .A1(_05420_),
    .S(_05603_),
    .X(_02333_));
 sky130_fd_sc_hd__mux2_1 _10589_ (.A0(\data_array.data1[1][1] ),
    .A1(_05422_),
    .S(_05603_),
    .X(_02334_));
 sky130_fd_sc_hd__mux2_1 _10590_ (.A0(\data_array.data1[1][2] ),
    .A1(_05424_),
    .S(_05603_),
    .X(_02335_));
 sky130_fd_sc_hd__mux2_1 _10591_ (.A0(\data_array.data1[1][3] ),
    .A1(_05426_),
    .S(_05603_),
    .X(_02336_));
 sky130_fd_sc_hd__mux2_1 _10592_ (.A0(\data_array.data1[1][4] ),
    .A1(_05428_),
    .S(_05603_),
    .X(_02337_));
 sky130_fd_sc_hd__mux2_1 _10593_ (.A0(\data_array.data1[1][5] ),
    .A1(_05430_),
    .S(_05603_),
    .X(_02338_));
 sky130_fd_sc_hd__mux2_1 _10594_ (.A0(\data_array.data1[1][6] ),
    .A1(_05432_),
    .S(_05603_),
    .X(_02339_));
 sky130_fd_sc_hd__mux2_1 _10595_ (.A0(\data_array.data1[1][7] ),
    .A1(_05434_),
    .S(_05603_),
    .X(_02340_));
 sky130_fd_sc_hd__mux2_1 _10596_ (.A0(\data_array.data1[1][8] ),
    .A1(_05436_),
    .S(_05603_),
    .X(_02341_));
 sky130_fd_sc_hd__mux2_1 _10597_ (.A0(\data_array.data1[1][9] ),
    .A1(_05438_),
    .S(_05603_),
    .X(_02342_));
 sky130_fd_sc_hd__mux2_1 _10598_ (.A0(\data_array.data1[1][10] ),
    .A1(_05440_),
    .S(_05603_),
    .X(_02343_));
 sky130_fd_sc_hd__mux2_1 _10599_ (.A0(\data_array.data1[1][11] ),
    .A1(_05442_),
    .S(_05603_),
    .X(_02344_));
 sky130_fd_sc_hd__mux2_1 _10600_ (.A0(\data_array.data1[1][12] ),
    .A1(_05444_),
    .S(_05603_),
    .X(_02345_));
 sky130_fd_sc_hd__mux2_1 _10601_ (.A0(\data_array.data1[1][13] ),
    .A1(_05446_),
    .S(_05603_),
    .X(_02346_));
 sky130_fd_sc_hd__mux2_1 _10602_ (.A0(\data_array.data1[1][14] ),
    .A1(_05448_),
    .S(_05603_),
    .X(_02347_));
 sky130_fd_sc_hd__mux2_1 _10603_ (.A0(\data_array.data1[1][15] ),
    .A1(_05450_),
    .S(_05603_),
    .X(_02348_));
 sky130_fd_sc_hd__mux2_1 _10604_ (.A0(\data_array.data1[1][16] ),
    .A1(_05452_),
    .S(_05603_),
    .X(_02349_));
 sky130_fd_sc_hd__mux2_1 _10605_ (.A0(\data_array.data1[1][17] ),
    .A1(_05454_),
    .S(_05603_),
    .X(_02350_));
 sky130_fd_sc_hd__mux2_1 _10606_ (.A0(\data_array.data1[1][18] ),
    .A1(_05456_),
    .S(_05603_),
    .X(_02351_));
 sky130_fd_sc_hd__mux2_1 _10607_ (.A0(\data_array.data1[1][19] ),
    .A1(_05458_),
    .S(_05603_),
    .X(_02352_));
 sky130_fd_sc_hd__mux2_1 _10608_ (.A0(\data_array.data1[1][20] ),
    .A1(_05460_),
    .S(_05603_),
    .X(_02353_));
 sky130_fd_sc_hd__mux2_1 _10609_ (.A0(\data_array.data1[1][21] ),
    .A1(_05462_),
    .S(_05603_),
    .X(_02354_));
 sky130_fd_sc_hd__mux2_1 _10610_ (.A0(\data_array.data1[1][22] ),
    .A1(_05464_),
    .S(_05603_),
    .X(_02355_));
 sky130_fd_sc_hd__mux2_1 _10611_ (.A0(\data_array.data1[1][23] ),
    .A1(_05466_),
    .S(_05603_),
    .X(_02356_));
 sky130_fd_sc_hd__mux2_1 _10612_ (.A0(\data_array.data1[1][24] ),
    .A1(_05468_),
    .S(_05603_),
    .X(_02357_));
 sky130_fd_sc_hd__mux2_1 _10613_ (.A0(\data_array.data1[1][25] ),
    .A1(_05470_),
    .S(_05603_),
    .X(_02358_));
 sky130_fd_sc_hd__mux2_1 _10614_ (.A0(\data_array.data1[1][26] ),
    .A1(_05472_),
    .S(_05603_),
    .X(_02359_));
 sky130_fd_sc_hd__mux2_1 _10615_ (.A0(\data_array.data1[1][27] ),
    .A1(_05474_),
    .S(_05603_),
    .X(_02360_));
 sky130_fd_sc_hd__mux2_1 _10616_ (.A0(\data_array.data1[1][28] ),
    .A1(_05476_),
    .S(_05603_),
    .X(_02361_));
 sky130_fd_sc_hd__mux2_1 _10617_ (.A0(\data_array.data1[1][29] ),
    .A1(_05478_),
    .S(_05603_),
    .X(_02362_));
 sky130_fd_sc_hd__mux2_1 _10618_ (.A0(\data_array.data1[1][30] ),
    .A1(_05480_),
    .S(_05603_),
    .X(_02363_));
 sky130_fd_sc_hd__mux2_1 _10619_ (.A0(\data_array.data1[1][31] ),
    .A1(_05482_),
    .S(_05603_),
    .X(_02364_));
 sky130_fd_sc_hd__mux2_1 _10620_ (.A0(\data_array.data1[1][32] ),
    .A1(_05484_),
    .S(_05603_),
    .X(_02365_));
 sky130_fd_sc_hd__mux2_1 _10621_ (.A0(\data_array.data1[1][33] ),
    .A1(_05486_),
    .S(_05603_),
    .X(_02366_));
 sky130_fd_sc_hd__mux2_1 _10622_ (.A0(\data_array.data1[1][34] ),
    .A1(_05488_),
    .S(_05603_),
    .X(_02367_));
 sky130_fd_sc_hd__mux2_1 _10623_ (.A0(\data_array.data1[1][35] ),
    .A1(_05490_),
    .S(_05603_),
    .X(_02368_));
 sky130_fd_sc_hd__mux2_1 _10624_ (.A0(\data_array.data1[1][36] ),
    .A1(_05492_),
    .S(_05603_),
    .X(_02369_));
 sky130_fd_sc_hd__mux2_1 _10625_ (.A0(\data_array.data1[1][37] ),
    .A1(_05494_),
    .S(_05603_),
    .X(_02370_));
 sky130_fd_sc_hd__mux2_1 _10626_ (.A0(\data_array.data1[1][38] ),
    .A1(_05496_),
    .S(_05603_),
    .X(_02371_));
 sky130_fd_sc_hd__mux2_1 _10627_ (.A0(\data_array.data1[1][39] ),
    .A1(_05498_),
    .S(_05603_),
    .X(_02372_));
 sky130_fd_sc_hd__mux2_1 _10628_ (.A0(\data_array.data1[1][40] ),
    .A1(_05500_),
    .S(_05603_),
    .X(_02373_));
 sky130_fd_sc_hd__mux2_1 _10629_ (.A0(\data_array.data1[1][41] ),
    .A1(_05502_),
    .S(_05603_),
    .X(_02374_));
 sky130_fd_sc_hd__mux2_1 _10630_ (.A0(\data_array.data1[1][42] ),
    .A1(_05504_),
    .S(_05603_),
    .X(_02375_));
 sky130_fd_sc_hd__mux2_1 _10631_ (.A0(\data_array.data1[1][43] ),
    .A1(_05506_),
    .S(_05603_),
    .X(_02376_));
 sky130_fd_sc_hd__mux2_1 _10632_ (.A0(\data_array.data1[1][44] ),
    .A1(_05508_),
    .S(_05603_),
    .X(_02377_));
 sky130_fd_sc_hd__mux2_1 _10633_ (.A0(\data_array.data1[1][45] ),
    .A1(_05510_),
    .S(_05603_),
    .X(_02378_));
 sky130_fd_sc_hd__mux2_1 _10634_ (.A0(\data_array.data1[1][46] ),
    .A1(_05512_),
    .S(_05603_),
    .X(_02379_));
 sky130_fd_sc_hd__mux2_1 _10635_ (.A0(\data_array.data1[1][47] ),
    .A1(_05514_),
    .S(_05603_),
    .X(_02380_));
 sky130_fd_sc_hd__mux2_1 _10636_ (.A0(\data_array.data1[1][48] ),
    .A1(_05516_),
    .S(_05603_),
    .X(_02381_));
 sky130_fd_sc_hd__mux2_1 _10637_ (.A0(\data_array.data1[1][49] ),
    .A1(_05518_),
    .S(_05603_),
    .X(_02382_));
 sky130_fd_sc_hd__mux2_1 _10638_ (.A0(\data_array.data1[1][50] ),
    .A1(_05520_),
    .S(_05603_),
    .X(_02383_));
 sky130_fd_sc_hd__mux2_1 _10639_ (.A0(\data_array.data1[1][51] ),
    .A1(_05522_),
    .S(_05603_),
    .X(_02384_));
 sky130_fd_sc_hd__mux2_1 _10640_ (.A0(\data_array.data1[1][52] ),
    .A1(_05524_),
    .S(_05603_),
    .X(_02385_));
 sky130_fd_sc_hd__mux2_1 _10641_ (.A0(\data_array.data1[1][53] ),
    .A1(_05526_),
    .S(_05603_),
    .X(_02386_));
 sky130_fd_sc_hd__mux2_1 _10642_ (.A0(\data_array.data1[1][54] ),
    .A1(_05528_),
    .S(_05603_),
    .X(_02387_));
 sky130_fd_sc_hd__mux2_1 _10643_ (.A0(\data_array.data1[1][55] ),
    .A1(_05530_),
    .S(_05603_),
    .X(_02388_));
 sky130_fd_sc_hd__mux2_1 _10644_ (.A0(\data_array.data1[1][56] ),
    .A1(_05532_),
    .S(_05603_),
    .X(_02389_));
 sky130_fd_sc_hd__mux2_1 _10645_ (.A0(\data_array.data1[1][57] ),
    .A1(_05534_),
    .S(_05603_),
    .X(_02390_));
 sky130_fd_sc_hd__mux2_1 _10646_ (.A0(\data_array.data1[1][58] ),
    .A1(_05536_),
    .S(_05603_),
    .X(_02391_));
 sky130_fd_sc_hd__mux2_1 _10647_ (.A0(\data_array.data1[1][59] ),
    .A1(_05538_),
    .S(_05603_),
    .X(_02392_));
 sky130_fd_sc_hd__mux2_1 _10648_ (.A0(\data_array.data1[1][60] ),
    .A1(_05540_),
    .S(_05603_),
    .X(_02393_));
 sky130_fd_sc_hd__mux2_1 _10649_ (.A0(\data_array.data1[1][61] ),
    .A1(_05542_),
    .S(_05603_),
    .X(_02394_));
 sky130_fd_sc_hd__mux2_1 _10650_ (.A0(\data_array.data1[1][62] ),
    .A1(_05544_),
    .S(_05603_),
    .X(_02395_));
 sky130_fd_sc_hd__mux2_1 _10651_ (.A0(\data_array.data1[1][63] ),
    .A1(_05546_),
    .S(_05603_),
    .X(_02396_));
 sky130_fd_sc_hd__mux2_1 _10652_ (.A0(\data_array.data1[2][0] ),
    .A1(_05420_),
    .S(_05602_),
    .X(_02397_));
 sky130_fd_sc_hd__mux2_1 _10653_ (.A0(\data_array.data1[2][1] ),
    .A1(_05422_),
    .S(_05602_),
    .X(_02398_));
 sky130_fd_sc_hd__mux2_1 _10654_ (.A0(\data_array.data1[2][2] ),
    .A1(_05424_),
    .S(_05602_),
    .X(_02399_));
 sky130_fd_sc_hd__mux2_1 _10655_ (.A0(\data_array.data1[2][3] ),
    .A1(_05426_),
    .S(_05602_),
    .X(_02400_));
 sky130_fd_sc_hd__mux2_1 _10656_ (.A0(\data_array.data1[2][4] ),
    .A1(_05428_),
    .S(_05602_),
    .X(_02401_));
 sky130_fd_sc_hd__mux2_1 _10657_ (.A0(\data_array.data1[2][5] ),
    .A1(_05430_),
    .S(_05602_),
    .X(_02402_));
 sky130_fd_sc_hd__mux2_1 _10658_ (.A0(\data_array.data1[2][6] ),
    .A1(_05432_),
    .S(_05602_),
    .X(_02403_));
 sky130_fd_sc_hd__mux2_1 _10659_ (.A0(\data_array.data1[2][7] ),
    .A1(_05434_),
    .S(_05602_),
    .X(_02404_));
 sky130_fd_sc_hd__mux2_1 _10660_ (.A0(\data_array.data1[2][8] ),
    .A1(_05436_),
    .S(_05602_),
    .X(_02405_));
 sky130_fd_sc_hd__mux2_1 _10661_ (.A0(\data_array.data1[2][9] ),
    .A1(_05438_),
    .S(_05602_),
    .X(_02406_));
 sky130_fd_sc_hd__mux2_1 _10662_ (.A0(\data_array.data1[2][10] ),
    .A1(_05440_),
    .S(_05602_),
    .X(_02407_));
 sky130_fd_sc_hd__mux2_1 _10663_ (.A0(\data_array.data1[2][11] ),
    .A1(_05442_),
    .S(_05602_),
    .X(_02408_));
 sky130_fd_sc_hd__mux2_1 _10664_ (.A0(\data_array.data1[2][12] ),
    .A1(_05444_),
    .S(_05602_),
    .X(_02409_));
 sky130_fd_sc_hd__mux2_1 _10665_ (.A0(\data_array.data1[2][13] ),
    .A1(_05446_),
    .S(_05602_),
    .X(_02410_));
 sky130_fd_sc_hd__mux2_1 _10666_ (.A0(\data_array.data1[2][14] ),
    .A1(_05448_),
    .S(_05602_),
    .X(_02411_));
 sky130_fd_sc_hd__mux2_1 _10667_ (.A0(\data_array.data1[2][15] ),
    .A1(_05450_),
    .S(_05602_),
    .X(_02412_));
 sky130_fd_sc_hd__mux2_1 _10668_ (.A0(\data_array.data1[2][16] ),
    .A1(_05452_),
    .S(_05602_),
    .X(_02413_));
 sky130_fd_sc_hd__mux2_1 _10669_ (.A0(\data_array.data1[2][17] ),
    .A1(_05454_),
    .S(_05602_),
    .X(_02414_));
 sky130_fd_sc_hd__mux2_1 _10670_ (.A0(\data_array.data1[2][18] ),
    .A1(_05456_),
    .S(_05602_),
    .X(_02415_));
 sky130_fd_sc_hd__mux2_1 _10671_ (.A0(\data_array.data1[2][19] ),
    .A1(_05458_),
    .S(_05602_),
    .X(_02416_));
 sky130_fd_sc_hd__mux2_1 _10672_ (.A0(\data_array.data1[2][20] ),
    .A1(_05460_),
    .S(_05602_),
    .X(_02417_));
 sky130_fd_sc_hd__mux2_1 _10673_ (.A0(\data_array.data1[2][21] ),
    .A1(_05462_),
    .S(_05602_),
    .X(_02418_));
 sky130_fd_sc_hd__mux2_1 _10674_ (.A0(\data_array.data1[2][22] ),
    .A1(_05464_),
    .S(_05602_),
    .X(_02419_));
 sky130_fd_sc_hd__mux2_1 _10675_ (.A0(\data_array.data1[2][23] ),
    .A1(_05466_),
    .S(_05602_),
    .X(_02420_));
 sky130_fd_sc_hd__mux2_1 _10676_ (.A0(\data_array.data1[2][24] ),
    .A1(_05468_),
    .S(_05602_),
    .X(_02421_));
 sky130_fd_sc_hd__mux2_1 _10677_ (.A0(\data_array.data1[2][25] ),
    .A1(_05470_),
    .S(_05602_),
    .X(_02422_));
 sky130_fd_sc_hd__mux2_1 _10678_ (.A0(\data_array.data1[2][26] ),
    .A1(_05472_),
    .S(_05602_),
    .X(_02423_));
 sky130_fd_sc_hd__mux2_1 _10679_ (.A0(\data_array.data1[2][27] ),
    .A1(_05474_),
    .S(_05602_),
    .X(_02424_));
 sky130_fd_sc_hd__mux2_1 _10680_ (.A0(\data_array.data1[2][28] ),
    .A1(_05476_),
    .S(_05602_),
    .X(_02425_));
 sky130_fd_sc_hd__mux2_1 _10681_ (.A0(\data_array.data1[2][29] ),
    .A1(_05478_),
    .S(_05602_),
    .X(_02426_));
 sky130_fd_sc_hd__mux2_1 _10682_ (.A0(\data_array.data1[2][30] ),
    .A1(_05480_),
    .S(_05602_),
    .X(_02427_));
 sky130_fd_sc_hd__mux2_1 _10683_ (.A0(\data_array.data1[2][31] ),
    .A1(_05482_),
    .S(_05602_),
    .X(_02428_));
 sky130_fd_sc_hd__mux2_1 _10684_ (.A0(\data_array.data1[2][32] ),
    .A1(_05484_),
    .S(_05602_),
    .X(_02429_));
 sky130_fd_sc_hd__mux2_1 _10685_ (.A0(\data_array.data1[2][33] ),
    .A1(_05486_),
    .S(_05602_),
    .X(_02430_));
 sky130_fd_sc_hd__mux2_1 _10686_ (.A0(\data_array.data1[2][34] ),
    .A1(_05488_),
    .S(_05602_),
    .X(_02431_));
 sky130_fd_sc_hd__mux2_1 _10687_ (.A0(\data_array.data1[2][35] ),
    .A1(_05490_),
    .S(_05602_),
    .X(_02432_));
 sky130_fd_sc_hd__mux2_1 _10688_ (.A0(\data_array.data1[2][36] ),
    .A1(_05492_),
    .S(_05602_),
    .X(_02433_));
 sky130_fd_sc_hd__mux2_1 _10689_ (.A0(\data_array.data1[2][37] ),
    .A1(_05494_),
    .S(_05602_),
    .X(_02434_));
 sky130_fd_sc_hd__mux2_1 _10690_ (.A0(\data_array.data1[2][38] ),
    .A1(_05496_),
    .S(_05602_),
    .X(_02435_));
 sky130_fd_sc_hd__mux2_1 _10691_ (.A0(\data_array.data1[2][39] ),
    .A1(_05498_),
    .S(_05602_),
    .X(_02436_));
 sky130_fd_sc_hd__mux2_1 _10692_ (.A0(\data_array.data1[2][40] ),
    .A1(_05500_),
    .S(_05602_),
    .X(_02437_));
 sky130_fd_sc_hd__mux2_1 _10693_ (.A0(\data_array.data1[2][41] ),
    .A1(_05502_),
    .S(_05602_),
    .X(_02438_));
 sky130_fd_sc_hd__mux2_1 _10694_ (.A0(\data_array.data1[2][42] ),
    .A1(_05504_),
    .S(_05602_),
    .X(_02439_));
 sky130_fd_sc_hd__mux2_1 _10695_ (.A0(\data_array.data1[2][43] ),
    .A1(_05506_),
    .S(_05602_),
    .X(_02440_));
 sky130_fd_sc_hd__mux2_1 _10696_ (.A0(\data_array.data1[2][44] ),
    .A1(_05508_),
    .S(_05602_),
    .X(_02441_));
 sky130_fd_sc_hd__mux2_1 _10697_ (.A0(\data_array.data1[2][45] ),
    .A1(_05510_),
    .S(_05602_),
    .X(_02442_));
 sky130_fd_sc_hd__mux2_1 _10698_ (.A0(\data_array.data1[2][46] ),
    .A1(_05512_),
    .S(_05602_),
    .X(_02443_));
 sky130_fd_sc_hd__mux2_1 _10699_ (.A0(\data_array.data1[2][47] ),
    .A1(_05514_),
    .S(_05602_),
    .X(_02444_));
 sky130_fd_sc_hd__mux2_1 _10700_ (.A0(\data_array.data1[2][48] ),
    .A1(_05516_),
    .S(_05602_),
    .X(_02445_));
 sky130_fd_sc_hd__mux2_1 _10701_ (.A0(\data_array.data1[2][49] ),
    .A1(_05518_),
    .S(_05602_),
    .X(_02446_));
 sky130_fd_sc_hd__mux2_1 _10702_ (.A0(\data_array.data1[2][50] ),
    .A1(_05520_),
    .S(_05602_),
    .X(_02447_));
 sky130_fd_sc_hd__mux2_1 _10703_ (.A0(\data_array.data1[2][51] ),
    .A1(_05522_),
    .S(_05602_),
    .X(_02448_));
 sky130_fd_sc_hd__mux2_1 _10704_ (.A0(\data_array.data1[2][52] ),
    .A1(_05524_),
    .S(_05602_),
    .X(_02449_));
 sky130_fd_sc_hd__mux2_1 _10705_ (.A0(\data_array.data1[2][53] ),
    .A1(_05526_),
    .S(_05602_),
    .X(_02450_));
 sky130_fd_sc_hd__mux2_1 _10706_ (.A0(\data_array.data1[2][54] ),
    .A1(_05528_),
    .S(_05602_),
    .X(_02451_));
 sky130_fd_sc_hd__mux2_1 _10707_ (.A0(\data_array.data1[2][55] ),
    .A1(_05530_),
    .S(_05602_),
    .X(_02452_));
 sky130_fd_sc_hd__mux2_1 _10708_ (.A0(\data_array.data1[2][56] ),
    .A1(_05532_),
    .S(_05602_),
    .X(_02453_));
 sky130_fd_sc_hd__mux2_1 _10709_ (.A0(\data_array.data1[2][57] ),
    .A1(_05534_),
    .S(_05602_),
    .X(_02454_));
 sky130_fd_sc_hd__mux2_1 _10710_ (.A0(\data_array.data1[2][58] ),
    .A1(_05536_),
    .S(_05602_),
    .X(_02455_));
 sky130_fd_sc_hd__mux2_1 _10711_ (.A0(\data_array.data1[2][59] ),
    .A1(_05538_),
    .S(_05602_),
    .X(_02456_));
 sky130_fd_sc_hd__mux2_1 _10712_ (.A0(\data_array.data1[2][60] ),
    .A1(_05540_),
    .S(_05602_),
    .X(_02457_));
 sky130_fd_sc_hd__mux2_1 _10713_ (.A0(\data_array.data1[2][61] ),
    .A1(_05542_),
    .S(_05602_),
    .X(_02458_));
 sky130_fd_sc_hd__mux2_1 _10714_ (.A0(\data_array.data1[2][62] ),
    .A1(_05544_),
    .S(_05602_),
    .X(_02459_));
 sky130_fd_sc_hd__mux2_1 _10715_ (.A0(\data_array.data1[2][63] ),
    .A1(_05546_),
    .S(_05602_),
    .X(_02460_));
 sky130_fd_sc_hd__mux2_1 _10716_ (.A0(_05420_),
    .A1(\data_array.data1[3][0] ),
    .S(_05601_),
    .X(_02461_));
 sky130_fd_sc_hd__mux2_1 _10717_ (.A0(_05422_),
    .A1(\data_array.data1[3][1] ),
    .S(_05601_),
    .X(_02462_));
 sky130_fd_sc_hd__mux2_1 _10718_ (.A0(_05424_),
    .A1(\data_array.data1[3][2] ),
    .S(_05601_),
    .X(_02463_));
 sky130_fd_sc_hd__mux2_1 _10719_ (.A0(_05426_),
    .A1(\data_array.data1[3][3] ),
    .S(_05601_),
    .X(_02464_));
 sky130_fd_sc_hd__mux2_1 _10720_ (.A0(_05428_),
    .A1(\data_array.data1[3][4] ),
    .S(_05601_),
    .X(_02465_));
 sky130_fd_sc_hd__mux2_1 _10721_ (.A0(_05430_),
    .A1(\data_array.data1[3][5] ),
    .S(_05601_),
    .X(_02466_));
 sky130_fd_sc_hd__mux2_1 _10722_ (.A0(_05432_),
    .A1(\data_array.data1[3][6] ),
    .S(_05601_),
    .X(_02467_));
 sky130_fd_sc_hd__mux2_1 _10723_ (.A0(_05434_),
    .A1(\data_array.data1[3][7] ),
    .S(_05601_),
    .X(_02468_));
 sky130_fd_sc_hd__mux2_1 _10724_ (.A0(_05436_),
    .A1(\data_array.data1[3][8] ),
    .S(_05601_),
    .X(_02469_));
 sky130_fd_sc_hd__mux2_1 _10725_ (.A0(_05438_),
    .A1(\data_array.data1[3][9] ),
    .S(_05601_),
    .X(_02470_));
 sky130_fd_sc_hd__mux2_1 _10726_ (.A0(_05440_),
    .A1(\data_array.data1[3][10] ),
    .S(_05601_),
    .X(_02471_));
 sky130_fd_sc_hd__mux2_1 _10727_ (.A0(_05442_),
    .A1(\data_array.data1[3][11] ),
    .S(_05601_),
    .X(_02472_));
 sky130_fd_sc_hd__mux2_1 _10728_ (.A0(_05444_),
    .A1(\data_array.data1[3][12] ),
    .S(_05601_),
    .X(_02473_));
 sky130_fd_sc_hd__mux2_1 _10729_ (.A0(_05446_),
    .A1(\data_array.data1[3][13] ),
    .S(_05601_),
    .X(_02474_));
 sky130_fd_sc_hd__mux2_1 _10730_ (.A0(_05448_),
    .A1(\data_array.data1[3][14] ),
    .S(_05601_),
    .X(_02475_));
 sky130_fd_sc_hd__mux2_1 _10731_ (.A0(_05450_),
    .A1(\data_array.data1[3][15] ),
    .S(_05601_),
    .X(_02476_));
 sky130_fd_sc_hd__mux2_1 _10732_ (.A0(_05452_),
    .A1(\data_array.data1[3][16] ),
    .S(_05601_),
    .X(_02477_));
 sky130_fd_sc_hd__mux2_1 _10733_ (.A0(_05454_),
    .A1(\data_array.data1[3][17] ),
    .S(_05601_),
    .X(_02478_));
 sky130_fd_sc_hd__mux2_1 _10734_ (.A0(_05456_),
    .A1(\data_array.data1[3][18] ),
    .S(_05601_),
    .X(_02479_));
 sky130_fd_sc_hd__mux2_1 _10735_ (.A0(_05458_),
    .A1(\data_array.data1[3][19] ),
    .S(_05601_),
    .X(_02480_));
 sky130_fd_sc_hd__mux2_1 _10736_ (.A0(_05460_),
    .A1(\data_array.data1[3][20] ),
    .S(_05601_),
    .X(_02481_));
 sky130_fd_sc_hd__mux2_1 _10737_ (.A0(_05462_),
    .A1(\data_array.data1[3][21] ),
    .S(_05601_),
    .X(_02482_));
 sky130_fd_sc_hd__mux2_1 _10738_ (.A0(_05464_),
    .A1(\data_array.data1[3][22] ),
    .S(_05601_),
    .X(_02483_));
 sky130_fd_sc_hd__mux2_1 _10739_ (.A0(_05466_),
    .A1(\data_array.data1[3][23] ),
    .S(_05601_),
    .X(_02484_));
 sky130_fd_sc_hd__mux2_1 _10740_ (.A0(_05468_),
    .A1(\data_array.data1[3][24] ),
    .S(_05601_),
    .X(_02485_));
 sky130_fd_sc_hd__mux2_1 _10741_ (.A0(_05470_),
    .A1(\data_array.data1[3][25] ),
    .S(_05601_),
    .X(_02486_));
 sky130_fd_sc_hd__mux2_1 _10742_ (.A0(_05472_),
    .A1(\data_array.data1[3][26] ),
    .S(_05601_),
    .X(_02487_));
 sky130_fd_sc_hd__mux2_1 _10743_ (.A0(_05474_),
    .A1(\data_array.data1[3][27] ),
    .S(_05601_),
    .X(_02488_));
 sky130_fd_sc_hd__mux2_1 _10744_ (.A0(_05476_),
    .A1(\data_array.data1[3][28] ),
    .S(_05601_),
    .X(_02489_));
 sky130_fd_sc_hd__mux2_1 _10745_ (.A0(_05478_),
    .A1(\data_array.data1[3][29] ),
    .S(_05601_),
    .X(_02490_));
 sky130_fd_sc_hd__mux2_1 _10746_ (.A0(_05480_),
    .A1(\data_array.data1[3][30] ),
    .S(_05601_),
    .X(_02491_));
 sky130_fd_sc_hd__mux2_1 _10747_ (.A0(_05482_),
    .A1(\data_array.data1[3][31] ),
    .S(_05601_),
    .X(_02492_));
 sky130_fd_sc_hd__mux2_1 _10748_ (.A0(_05484_),
    .A1(\data_array.data1[3][32] ),
    .S(_05601_),
    .X(_02493_));
 sky130_fd_sc_hd__mux2_1 _10749_ (.A0(_05486_),
    .A1(\data_array.data1[3][33] ),
    .S(_05601_),
    .X(_02494_));
 sky130_fd_sc_hd__mux2_1 _10750_ (.A0(_05488_),
    .A1(\data_array.data1[3][34] ),
    .S(_05601_),
    .X(_02495_));
 sky130_fd_sc_hd__mux2_1 _10751_ (.A0(_05490_),
    .A1(\data_array.data1[3][35] ),
    .S(_05601_),
    .X(_02496_));
 sky130_fd_sc_hd__mux2_1 _10752_ (.A0(_05492_),
    .A1(\data_array.data1[3][36] ),
    .S(_05601_),
    .X(_02497_));
 sky130_fd_sc_hd__mux2_1 _10753_ (.A0(_05494_),
    .A1(\data_array.data1[3][37] ),
    .S(_05601_),
    .X(_02498_));
 sky130_fd_sc_hd__mux2_1 _10754_ (.A0(_05496_),
    .A1(\data_array.data1[3][38] ),
    .S(_05601_),
    .X(_02499_));
 sky130_fd_sc_hd__mux2_1 _10755_ (.A0(_05498_),
    .A1(\data_array.data1[3][39] ),
    .S(_05601_),
    .X(_02500_));
 sky130_fd_sc_hd__mux2_1 _10756_ (.A0(_05500_),
    .A1(\data_array.data1[3][40] ),
    .S(_05601_),
    .X(_02501_));
 sky130_fd_sc_hd__mux2_1 _10757_ (.A0(_05502_),
    .A1(\data_array.data1[3][41] ),
    .S(_05601_),
    .X(_02502_));
 sky130_fd_sc_hd__mux2_1 _10758_ (.A0(_05504_),
    .A1(\data_array.data1[3][42] ),
    .S(_05601_),
    .X(_02503_));
 sky130_fd_sc_hd__mux2_1 _10759_ (.A0(_05506_),
    .A1(\data_array.data1[3][43] ),
    .S(_05601_),
    .X(_02504_));
 sky130_fd_sc_hd__mux2_1 _10760_ (.A0(_05508_),
    .A1(\data_array.data1[3][44] ),
    .S(_05601_),
    .X(_02505_));
 sky130_fd_sc_hd__mux2_1 _10761_ (.A0(_05510_),
    .A1(\data_array.data1[3][45] ),
    .S(_05601_),
    .X(_02506_));
 sky130_fd_sc_hd__mux2_1 _10762_ (.A0(_05512_),
    .A1(\data_array.data1[3][46] ),
    .S(_05601_),
    .X(_02507_));
 sky130_fd_sc_hd__mux2_1 _10763_ (.A0(_05514_),
    .A1(\data_array.data1[3][47] ),
    .S(_05601_),
    .X(_02508_));
 sky130_fd_sc_hd__mux2_1 _10764_ (.A0(_05516_),
    .A1(\data_array.data1[3][48] ),
    .S(_05601_),
    .X(_02509_));
 sky130_fd_sc_hd__mux2_1 _10765_ (.A0(_05518_),
    .A1(\data_array.data1[3][49] ),
    .S(_05601_),
    .X(_02510_));
 sky130_fd_sc_hd__mux2_1 _10766_ (.A0(_05520_),
    .A1(\data_array.data1[3][50] ),
    .S(_05601_),
    .X(_02511_));
 sky130_fd_sc_hd__mux2_1 _10767_ (.A0(_05522_),
    .A1(\data_array.data1[3][51] ),
    .S(_05601_),
    .X(_02512_));
 sky130_fd_sc_hd__mux2_1 _10768_ (.A0(_05524_),
    .A1(\data_array.data1[3][52] ),
    .S(_05601_),
    .X(_02513_));
 sky130_fd_sc_hd__mux2_1 _10769_ (.A0(_05526_),
    .A1(\data_array.data1[3][53] ),
    .S(_05601_),
    .X(_02514_));
 sky130_fd_sc_hd__mux2_1 _10770_ (.A0(_05528_),
    .A1(\data_array.data1[3][54] ),
    .S(_05601_),
    .X(_02515_));
 sky130_fd_sc_hd__mux2_1 _10771_ (.A0(_05530_),
    .A1(\data_array.data1[3][55] ),
    .S(_05601_),
    .X(_02516_));
 sky130_fd_sc_hd__mux2_1 _10772_ (.A0(_05532_),
    .A1(\data_array.data1[3][56] ),
    .S(_05601_),
    .X(_02517_));
 sky130_fd_sc_hd__mux2_1 _10773_ (.A0(_05534_),
    .A1(\data_array.data1[3][57] ),
    .S(_05601_),
    .X(_02518_));
 sky130_fd_sc_hd__mux2_1 _10774_ (.A0(_05536_),
    .A1(\data_array.data1[3][58] ),
    .S(_05601_),
    .X(_02519_));
 sky130_fd_sc_hd__mux2_1 _10775_ (.A0(_05538_),
    .A1(\data_array.data1[3][59] ),
    .S(_05601_),
    .X(_02520_));
 sky130_fd_sc_hd__mux2_1 _10776_ (.A0(_05540_),
    .A1(\data_array.data1[3][60] ),
    .S(_05601_),
    .X(_02521_));
 sky130_fd_sc_hd__mux2_1 _10777_ (.A0(_05542_),
    .A1(\data_array.data1[3][61] ),
    .S(_05601_),
    .X(_02522_));
 sky130_fd_sc_hd__mux2_1 _10778_ (.A0(_05544_),
    .A1(\data_array.data1[3][62] ),
    .S(_05601_),
    .X(_02523_));
 sky130_fd_sc_hd__mux2_1 _10779_ (.A0(_05546_),
    .A1(\data_array.data1[3][63] ),
    .S(_05601_),
    .X(_02524_));
 sky130_fd_sc_hd__mux2_1 _10780_ (.A0(\data_array.data1[4][0] ),
    .A1(_05420_),
    .S(_05600_),
    .X(_02525_));
 sky130_fd_sc_hd__mux2_1 _10781_ (.A0(\data_array.data1[4][1] ),
    .A1(_05422_),
    .S(_05600_),
    .X(_02526_));
 sky130_fd_sc_hd__mux2_1 _10782_ (.A0(\data_array.data1[4][2] ),
    .A1(_05424_),
    .S(_05600_),
    .X(_02527_));
 sky130_fd_sc_hd__mux2_1 _10783_ (.A0(\data_array.data1[4][3] ),
    .A1(_05426_),
    .S(_05600_),
    .X(_02528_));
 sky130_fd_sc_hd__mux2_1 _10784_ (.A0(\data_array.data1[4][4] ),
    .A1(_05428_),
    .S(_05600_),
    .X(_02529_));
 sky130_fd_sc_hd__mux2_1 _10785_ (.A0(\data_array.data1[4][5] ),
    .A1(_05430_),
    .S(_05600_),
    .X(_02530_));
 sky130_fd_sc_hd__mux2_1 _10786_ (.A0(\data_array.data1[4][6] ),
    .A1(_05432_),
    .S(_05600_),
    .X(_02531_));
 sky130_fd_sc_hd__mux2_1 _10787_ (.A0(\data_array.data1[4][7] ),
    .A1(_05434_),
    .S(_05600_),
    .X(_02532_));
 sky130_fd_sc_hd__mux2_1 _10788_ (.A0(\data_array.data1[4][8] ),
    .A1(_05436_),
    .S(_05600_),
    .X(_02533_));
 sky130_fd_sc_hd__mux2_1 _10789_ (.A0(\data_array.data1[4][9] ),
    .A1(_05438_),
    .S(_05600_),
    .X(_02534_));
 sky130_fd_sc_hd__mux2_1 _10790_ (.A0(\data_array.data1[4][10] ),
    .A1(_05440_),
    .S(_05600_),
    .X(_02535_));
 sky130_fd_sc_hd__mux2_1 _10791_ (.A0(\data_array.data1[4][11] ),
    .A1(_05442_),
    .S(_05600_),
    .X(_02536_));
 sky130_fd_sc_hd__mux2_1 _10792_ (.A0(\data_array.data1[4][12] ),
    .A1(_05444_),
    .S(_05600_),
    .X(_02537_));
 sky130_fd_sc_hd__mux2_1 _10793_ (.A0(\data_array.data1[4][13] ),
    .A1(_05446_),
    .S(_05600_),
    .X(_02538_));
 sky130_fd_sc_hd__mux2_1 _10794_ (.A0(\data_array.data1[4][14] ),
    .A1(_05448_),
    .S(_05600_),
    .X(_02539_));
 sky130_fd_sc_hd__mux2_1 _10795_ (.A0(\data_array.data1[4][15] ),
    .A1(_05450_),
    .S(_05600_),
    .X(_02540_));
 sky130_fd_sc_hd__mux2_1 _10796_ (.A0(\data_array.data1[4][16] ),
    .A1(_05452_),
    .S(_05600_),
    .X(_02541_));
 sky130_fd_sc_hd__mux2_1 _10797_ (.A0(\data_array.data1[4][17] ),
    .A1(_05454_),
    .S(_05600_),
    .X(_02542_));
 sky130_fd_sc_hd__mux2_1 _10798_ (.A0(\data_array.data1[4][18] ),
    .A1(_05456_),
    .S(_05600_),
    .X(_02543_));
 sky130_fd_sc_hd__mux2_1 _10799_ (.A0(\data_array.data1[4][19] ),
    .A1(_05458_),
    .S(_05600_),
    .X(_02544_));
 sky130_fd_sc_hd__mux2_1 _10800_ (.A0(\data_array.data1[4][20] ),
    .A1(_05460_),
    .S(_05600_),
    .X(_02545_));
 sky130_fd_sc_hd__mux2_1 _10801_ (.A0(\data_array.data1[4][21] ),
    .A1(_05462_),
    .S(_05600_),
    .X(_02546_));
 sky130_fd_sc_hd__mux2_1 _10802_ (.A0(\data_array.data1[4][22] ),
    .A1(_05464_),
    .S(_05600_),
    .X(_02547_));
 sky130_fd_sc_hd__mux2_1 _10803_ (.A0(\data_array.data1[4][23] ),
    .A1(_05466_),
    .S(_05600_),
    .X(_02548_));
 sky130_fd_sc_hd__mux2_1 _10804_ (.A0(\data_array.data1[4][24] ),
    .A1(_05468_),
    .S(_05600_),
    .X(_02549_));
 sky130_fd_sc_hd__mux2_1 _10805_ (.A0(\data_array.data1[4][25] ),
    .A1(_05470_),
    .S(_05600_),
    .X(_02550_));
 sky130_fd_sc_hd__mux2_1 _10806_ (.A0(\data_array.data1[4][26] ),
    .A1(_05472_),
    .S(_05600_),
    .X(_02551_));
 sky130_fd_sc_hd__mux2_1 _10807_ (.A0(\data_array.data1[4][27] ),
    .A1(_05474_),
    .S(_05600_),
    .X(_02552_));
 sky130_fd_sc_hd__mux2_1 _10808_ (.A0(\data_array.data1[4][28] ),
    .A1(_05476_),
    .S(_05600_),
    .X(_02553_));
 sky130_fd_sc_hd__mux2_1 _10809_ (.A0(\data_array.data1[4][29] ),
    .A1(_05478_),
    .S(_05600_),
    .X(_02554_));
 sky130_fd_sc_hd__mux2_1 _10810_ (.A0(\data_array.data1[4][30] ),
    .A1(_05480_),
    .S(_05600_),
    .X(_02555_));
 sky130_fd_sc_hd__mux2_1 _10811_ (.A0(\data_array.data1[4][31] ),
    .A1(_05482_),
    .S(_05600_),
    .X(_02556_));
 sky130_fd_sc_hd__mux2_1 _10812_ (.A0(\data_array.data1[4][32] ),
    .A1(_05484_),
    .S(_05600_),
    .X(_02557_));
 sky130_fd_sc_hd__mux2_1 _10813_ (.A0(\data_array.data1[4][33] ),
    .A1(_05486_),
    .S(_05600_),
    .X(_02558_));
 sky130_fd_sc_hd__mux2_1 _10814_ (.A0(\data_array.data1[4][34] ),
    .A1(_05488_),
    .S(_05600_),
    .X(_02559_));
 sky130_fd_sc_hd__mux2_1 _10815_ (.A0(\data_array.data1[4][35] ),
    .A1(_05490_),
    .S(_05600_),
    .X(_02560_));
 sky130_fd_sc_hd__mux2_1 _10816_ (.A0(\data_array.data1[4][36] ),
    .A1(_05492_),
    .S(_05600_),
    .X(_02561_));
 sky130_fd_sc_hd__mux2_1 _10817_ (.A0(\data_array.data1[4][37] ),
    .A1(_05494_),
    .S(_05600_),
    .X(_02562_));
 sky130_fd_sc_hd__mux2_1 _10818_ (.A0(\data_array.data1[4][38] ),
    .A1(_05496_),
    .S(_05600_),
    .X(_02563_));
 sky130_fd_sc_hd__mux2_1 _10819_ (.A0(\data_array.data1[4][39] ),
    .A1(_05498_),
    .S(_05600_),
    .X(_02564_));
 sky130_fd_sc_hd__mux2_1 _10820_ (.A0(\data_array.data1[4][40] ),
    .A1(_05500_),
    .S(_05600_),
    .X(_02565_));
 sky130_fd_sc_hd__mux2_1 _10821_ (.A0(\data_array.data1[4][41] ),
    .A1(_05502_),
    .S(_05600_),
    .X(_02566_));
 sky130_fd_sc_hd__mux2_1 _10822_ (.A0(\data_array.data1[4][42] ),
    .A1(_05504_),
    .S(_05600_),
    .X(_02567_));
 sky130_fd_sc_hd__mux2_1 _10823_ (.A0(\data_array.data1[4][43] ),
    .A1(_05506_),
    .S(_05600_),
    .X(_02568_));
 sky130_fd_sc_hd__mux2_1 _10824_ (.A0(\data_array.data1[4][44] ),
    .A1(_05508_),
    .S(_05600_),
    .X(_02569_));
 sky130_fd_sc_hd__mux2_1 _10825_ (.A0(\data_array.data1[4][45] ),
    .A1(_05510_),
    .S(_05600_),
    .X(_02570_));
 sky130_fd_sc_hd__mux2_1 _10826_ (.A0(\data_array.data1[4][46] ),
    .A1(_05512_),
    .S(_05600_),
    .X(_02571_));
 sky130_fd_sc_hd__mux2_1 _10827_ (.A0(\data_array.data1[4][47] ),
    .A1(_05514_),
    .S(_05600_),
    .X(_02572_));
 sky130_fd_sc_hd__mux2_1 _10828_ (.A0(\data_array.data1[4][48] ),
    .A1(_05516_),
    .S(_05600_),
    .X(_02573_));
 sky130_fd_sc_hd__mux2_1 _10829_ (.A0(\data_array.data1[4][49] ),
    .A1(_05518_),
    .S(_05600_),
    .X(_02574_));
 sky130_fd_sc_hd__mux2_1 _10830_ (.A0(\data_array.data1[4][50] ),
    .A1(_05520_),
    .S(_05600_),
    .X(_02575_));
 sky130_fd_sc_hd__mux2_1 _10831_ (.A0(\data_array.data1[4][51] ),
    .A1(_05522_),
    .S(_05600_),
    .X(_02576_));
 sky130_fd_sc_hd__mux2_1 _10832_ (.A0(\data_array.data1[4][52] ),
    .A1(_05524_),
    .S(_05600_),
    .X(_02577_));
 sky130_fd_sc_hd__mux2_1 _10833_ (.A0(\data_array.data1[4][53] ),
    .A1(_05526_),
    .S(_05600_),
    .X(_02578_));
 sky130_fd_sc_hd__mux2_1 _10834_ (.A0(\data_array.data1[4][54] ),
    .A1(_05528_),
    .S(_05600_),
    .X(_02579_));
 sky130_fd_sc_hd__mux2_1 _10835_ (.A0(\data_array.data1[4][55] ),
    .A1(_05530_),
    .S(_05600_),
    .X(_02580_));
 sky130_fd_sc_hd__mux2_1 _10836_ (.A0(\data_array.data1[4][56] ),
    .A1(_05532_),
    .S(_05600_),
    .X(_02581_));
 sky130_fd_sc_hd__mux2_1 _10837_ (.A0(\data_array.data1[4][57] ),
    .A1(_05534_),
    .S(_05600_),
    .X(_02582_));
 sky130_fd_sc_hd__mux2_1 _10838_ (.A0(\data_array.data1[4][58] ),
    .A1(_05536_),
    .S(_05600_),
    .X(_02583_));
 sky130_fd_sc_hd__mux2_1 _10839_ (.A0(\data_array.data1[4][59] ),
    .A1(_05538_),
    .S(_05600_),
    .X(_02584_));
 sky130_fd_sc_hd__mux2_1 _10840_ (.A0(\data_array.data1[4][60] ),
    .A1(_05540_),
    .S(_05600_),
    .X(_02585_));
 sky130_fd_sc_hd__mux2_1 _10841_ (.A0(\data_array.data1[4][61] ),
    .A1(_05542_),
    .S(_05600_),
    .X(_02586_));
 sky130_fd_sc_hd__mux2_1 _10842_ (.A0(\data_array.data1[4][62] ),
    .A1(_05544_),
    .S(_05600_),
    .X(_02587_));
 sky130_fd_sc_hd__mux2_1 _10843_ (.A0(\data_array.data1[4][63] ),
    .A1(_05546_),
    .S(_05600_),
    .X(_02588_));
 sky130_fd_sc_hd__mux2_1 _10844_ (.A0(_05420_),
    .A1(\data_array.data1[5][0] ),
    .S(_05599_),
    .X(_02589_));
 sky130_fd_sc_hd__mux2_1 _10845_ (.A0(_05422_),
    .A1(\data_array.data1[5][1] ),
    .S(_05599_),
    .X(_02590_));
 sky130_fd_sc_hd__mux2_1 _10846_ (.A0(_05424_),
    .A1(\data_array.data1[5][2] ),
    .S(_05599_),
    .X(_02591_));
 sky130_fd_sc_hd__mux2_1 _10847_ (.A0(_05426_),
    .A1(\data_array.data1[5][3] ),
    .S(_05599_),
    .X(_02592_));
 sky130_fd_sc_hd__mux2_1 _10848_ (.A0(_05428_),
    .A1(\data_array.data1[5][4] ),
    .S(_05599_),
    .X(_02593_));
 sky130_fd_sc_hd__mux2_1 _10849_ (.A0(_05430_),
    .A1(\data_array.data1[5][5] ),
    .S(_05599_),
    .X(_02594_));
 sky130_fd_sc_hd__mux2_1 _10850_ (.A0(_05432_),
    .A1(\data_array.data1[5][6] ),
    .S(_05599_),
    .X(_02595_));
 sky130_fd_sc_hd__mux2_1 _10851_ (.A0(_05434_),
    .A1(\data_array.data1[5][7] ),
    .S(_05599_),
    .X(_02596_));
 sky130_fd_sc_hd__mux2_1 _10852_ (.A0(_05436_),
    .A1(\data_array.data1[5][8] ),
    .S(_05599_),
    .X(_02597_));
 sky130_fd_sc_hd__mux2_1 _10853_ (.A0(_05438_),
    .A1(\data_array.data1[5][9] ),
    .S(_05599_),
    .X(_02598_));
 sky130_fd_sc_hd__mux2_1 _10854_ (.A0(_05440_),
    .A1(\data_array.data1[5][10] ),
    .S(_05599_),
    .X(_02599_));
 sky130_fd_sc_hd__mux2_1 _10855_ (.A0(_05442_),
    .A1(\data_array.data1[5][11] ),
    .S(_05599_),
    .X(_02600_));
 sky130_fd_sc_hd__mux2_1 _10856_ (.A0(_05444_),
    .A1(\data_array.data1[5][12] ),
    .S(_05599_),
    .X(_02601_));
 sky130_fd_sc_hd__mux2_1 _10857_ (.A0(_05446_),
    .A1(\data_array.data1[5][13] ),
    .S(_05599_),
    .X(_02602_));
 sky130_fd_sc_hd__mux2_1 _10858_ (.A0(_05448_),
    .A1(\data_array.data1[5][14] ),
    .S(_05599_),
    .X(_02603_));
 sky130_fd_sc_hd__mux2_1 _10859_ (.A0(_05450_),
    .A1(\data_array.data1[5][15] ),
    .S(_05599_),
    .X(_02604_));
 sky130_fd_sc_hd__mux2_1 _10860_ (.A0(_05452_),
    .A1(\data_array.data1[5][16] ),
    .S(_05599_),
    .X(_02605_));
 sky130_fd_sc_hd__mux2_1 _10861_ (.A0(_05454_),
    .A1(\data_array.data1[5][17] ),
    .S(_05599_),
    .X(_02606_));
 sky130_fd_sc_hd__mux2_1 _10862_ (.A0(_05456_),
    .A1(\data_array.data1[5][18] ),
    .S(_05599_),
    .X(_02607_));
 sky130_fd_sc_hd__mux2_1 _10863_ (.A0(_05458_),
    .A1(\data_array.data1[5][19] ),
    .S(_05599_),
    .X(_02608_));
 sky130_fd_sc_hd__mux2_1 _10864_ (.A0(_05460_),
    .A1(\data_array.data1[5][20] ),
    .S(_05599_),
    .X(_02609_));
 sky130_fd_sc_hd__mux2_1 _10865_ (.A0(_05462_),
    .A1(\data_array.data1[5][21] ),
    .S(_05599_),
    .X(_02610_));
 sky130_fd_sc_hd__mux2_1 _10866_ (.A0(_05464_),
    .A1(\data_array.data1[5][22] ),
    .S(_05599_),
    .X(_02611_));
 sky130_fd_sc_hd__mux2_1 _10867_ (.A0(_05466_),
    .A1(\data_array.data1[5][23] ),
    .S(_05599_),
    .X(_02612_));
 sky130_fd_sc_hd__mux2_1 _10868_ (.A0(_05468_),
    .A1(\data_array.data1[5][24] ),
    .S(_05599_),
    .X(_02613_));
 sky130_fd_sc_hd__mux2_1 _10869_ (.A0(_05470_),
    .A1(\data_array.data1[5][25] ),
    .S(_05599_),
    .X(_02614_));
 sky130_fd_sc_hd__mux2_1 _10870_ (.A0(_05472_),
    .A1(\data_array.data1[5][26] ),
    .S(_05599_),
    .X(_02615_));
 sky130_fd_sc_hd__mux2_1 _10871_ (.A0(_05474_),
    .A1(\data_array.data1[5][27] ),
    .S(_05599_),
    .X(_02616_));
 sky130_fd_sc_hd__mux2_1 _10872_ (.A0(_05476_),
    .A1(\data_array.data1[5][28] ),
    .S(_05599_),
    .X(_02617_));
 sky130_fd_sc_hd__mux2_1 _10873_ (.A0(_05478_),
    .A1(\data_array.data1[5][29] ),
    .S(_05599_),
    .X(_02618_));
 sky130_fd_sc_hd__mux2_1 _10874_ (.A0(_05480_),
    .A1(\data_array.data1[5][30] ),
    .S(_05599_),
    .X(_02619_));
 sky130_fd_sc_hd__mux2_1 _10875_ (.A0(_05482_),
    .A1(\data_array.data1[5][31] ),
    .S(_05599_),
    .X(_02620_));
 sky130_fd_sc_hd__mux2_1 _10876_ (.A0(_05484_),
    .A1(\data_array.data1[5][32] ),
    .S(_05599_),
    .X(_02621_));
 sky130_fd_sc_hd__mux2_1 _10877_ (.A0(_05486_),
    .A1(\data_array.data1[5][33] ),
    .S(_05599_),
    .X(_02622_));
 sky130_fd_sc_hd__mux2_1 _10878_ (.A0(_05488_),
    .A1(\data_array.data1[5][34] ),
    .S(_05599_),
    .X(_02623_));
 sky130_fd_sc_hd__mux2_1 _10879_ (.A0(_05490_),
    .A1(\data_array.data1[5][35] ),
    .S(_05599_),
    .X(_02624_));
 sky130_fd_sc_hd__mux2_1 _10880_ (.A0(_05492_),
    .A1(\data_array.data1[5][36] ),
    .S(_05599_),
    .X(_02625_));
 sky130_fd_sc_hd__mux2_1 _10881_ (.A0(_05494_),
    .A1(\data_array.data1[5][37] ),
    .S(_05599_),
    .X(_02626_));
 sky130_fd_sc_hd__mux2_1 _10882_ (.A0(_05496_),
    .A1(\data_array.data1[5][38] ),
    .S(_05599_),
    .X(_02627_));
 sky130_fd_sc_hd__mux2_1 _10883_ (.A0(_05498_),
    .A1(\data_array.data1[5][39] ),
    .S(_05599_),
    .X(_02628_));
 sky130_fd_sc_hd__mux2_1 _10884_ (.A0(_05500_),
    .A1(\data_array.data1[5][40] ),
    .S(_05599_),
    .X(_02629_));
 sky130_fd_sc_hd__mux2_1 _10885_ (.A0(_05502_),
    .A1(\data_array.data1[5][41] ),
    .S(_05599_),
    .X(_02630_));
 sky130_fd_sc_hd__mux2_1 _10886_ (.A0(_05504_),
    .A1(\data_array.data1[5][42] ),
    .S(_05599_),
    .X(_02631_));
 sky130_fd_sc_hd__mux2_1 _10887_ (.A0(_05506_),
    .A1(\data_array.data1[5][43] ),
    .S(_05599_),
    .X(_02632_));
 sky130_fd_sc_hd__mux2_1 _10888_ (.A0(_05508_),
    .A1(\data_array.data1[5][44] ),
    .S(_05599_),
    .X(_02633_));
 sky130_fd_sc_hd__mux2_1 _10889_ (.A0(_05510_),
    .A1(\data_array.data1[5][45] ),
    .S(_05599_),
    .X(_02634_));
 sky130_fd_sc_hd__mux2_1 _10890_ (.A0(_05512_),
    .A1(\data_array.data1[5][46] ),
    .S(_05599_),
    .X(_02635_));
 sky130_fd_sc_hd__mux2_1 _10891_ (.A0(_05514_),
    .A1(\data_array.data1[5][47] ),
    .S(_05599_),
    .X(_02636_));
 sky130_fd_sc_hd__mux2_1 _10892_ (.A0(_05516_),
    .A1(\data_array.data1[5][48] ),
    .S(_05599_),
    .X(_02637_));
 sky130_fd_sc_hd__mux2_1 _10893_ (.A0(_05518_),
    .A1(\data_array.data1[5][49] ),
    .S(_05599_),
    .X(_02638_));
 sky130_fd_sc_hd__mux2_1 _10894_ (.A0(_05520_),
    .A1(\data_array.data1[5][50] ),
    .S(_05599_),
    .X(_02639_));
 sky130_fd_sc_hd__mux2_1 _10895_ (.A0(_05522_),
    .A1(\data_array.data1[5][51] ),
    .S(_05599_),
    .X(_02640_));
 sky130_fd_sc_hd__mux2_1 _10896_ (.A0(_05524_),
    .A1(\data_array.data1[5][52] ),
    .S(_05599_),
    .X(_02641_));
 sky130_fd_sc_hd__mux2_1 _10897_ (.A0(_05526_),
    .A1(\data_array.data1[5][53] ),
    .S(_05599_),
    .X(_02642_));
 sky130_fd_sc_hd__mux2_1 _10898_ (.A0(_05528_),
    .A1(\data_array.data1[5][54] ),
    .S(_05599_),
    .X(_02643_));
 sky130_fd_sc_hd__mux2_1 _10899_ (.A0(_05530_),
    .A1(\data_array.data1[5][55] ),
    .S(_05599_),
    .X(_02644_));
 sky130_fd_sc_hd__mux2_1 _10900_ (.A0(_05532_),
    .A1(\data_array.data1[5][56] ),
    .S(_05599_),
    .X(_02645_));
 sky130_fd_sc_hd__mux2_1 _10901_ (.A0(_05534_),
    .A1(\data_array.data1[5][57] ),
    .S(_05599_),
    .X(_02646_));
 sky130_fd_sc_hd__mux2_1 _10902_ (.A0(_05536_),
    .A1(\data_array.data1[5][58] ),
    .S(_05599_),
    .X(_02647_));
 sky130_fd_sc_hd__mux2_1 _10903_ (.A0(_05538_),
    .A1(\data_array.data1[5][59] ),
    .S(_05599_),
    .X(_02648_));
 sky130_fd_sc_hd__mux2_1 _10904_ (.A0(_05540_),
    .A1(\data_array.data1[5][60] ),
    .S(_05599_),
    .X(_02649_));
 sky130_fd_sc_hd__mux2_1 _10905_ (.A0(_05542_),
    .A1(\data_array.data1[5][61] ),
    .S(_05599_),
    .X(_02650_));
 sky130_fd_sc_hd__mux2_1 _10906_ (.A0(_05544_),
    .A1(\data_array.data1[5][62] ),
    .S(_05599_),
    .X(_02651_));
 sky130_fd_sc_hd__mux2_1 _10907_ (.A0(_05546_),
    .A1(\data_array.data1[5][63] ),
    .S(_05599_),
    .X(_02652_));
 sky130_fd_sc_hd__mux2_1 _10908_ (.A0(_05420_),
    .A1(\data_array.data1[6][0] ),
    .S(_05598_),
    .X(_02653_));
 sky130_fd_sc_hd__mux2_1 _10909_ (.A0(_05422_),
    .A1(\data_array.data1[6][1] ),
    .S(_05598_),
    .X(_02654_));
 sky130_fd_sc_hd__mux2_1 _10910_ (.A0(_05424_),
    .A1(\data_array.data1[6][2] ),
    .S(_05598_),
    .X(_02655_));
 sky130_fd_sc_hd__mux2_1 _10911_ (.A0(_05426_),
    .A1(\data_array.data1[6][3] ),
    .S(_05598_),
    .X(_02656_));
 sky130_fd_sc_hd__mux2_1 _10912_ (.A0(_05428_),
    .A1(\data_array.data1[6][4] ),
    .S(_05598_),
    .X(_02657_));
 sky130_fd_sc_hd__mux2_1 _10913_ (.A0(_05430_),
    .A1(\data_array.data1[6][5] ),
    .S(_05598_),
    .X(_02658_));
 sky130_fd_sc_hd__mux2_1 _10914_ (.A0(_05432_),
    .A1(\data_array.data1[6][6] ),
    .S(_05598_),
    .X(_02659_));
 sky130_fd_sc_hd__mux2_1 _10915_ (.A0(_05434_),
    .A1(\data_array.data1[6][7] ),
    .S(_05598_),
    .X(_02660_));
 sky130_fd_sc_hd__mux2_1 _10916_ (.A0(_05436_),
    .A1(\data_array.data1[6][8] ),
    .S(_05598_),
    .X(_02661_));
 sky130_fd_sc_hd__mux2_1 _10917_ (.A0(_05438_),
    .A1(\data_array.data1[6][9] ),
    .S(_05598_),
    .X(_02662_));
 sky130_fd_sc_hd__mux2_1 _10918_ (.A0(_05440_),
    .A1(\data_array.data1[6][10] ),
    .S(_05598_),
    .X(_02663_));
 sky130_fd_sc_hd__mux2_1 _10919_ (.A0(_05442_),
    .A1(\data_array.data1[6][11] ),
    .S(_05598_),
    .X(_02664_));
 sky130_fd_sc_hd__mux2_1 _10920_ (.A0(_05444_),
    .A1(\data_array.data1[6][12] ),
    .S(_05598_),
    .X(_02665_));
 sky130_fd_sc_hd__mux2_1 _10921_ (.A0(_05446_),
    .A1(\data_array.data1[6][13] ),
    .S(_05598_),
    .X(_02666_));
 sky130_fd_sc_hd__mux2_1 _10922_ (.A0(_05448_),
    .A1(\data_array.data1[6][14] ),
    .S(_05598_),
    .X(_02667_));
 sky130_fd_sc_hd__mux2_1 _10923_ (.A0(_05450_),
    .A1(\data_array.data1[6][15] ),
    .S(_05598_),
    .X(_02668_));
 sky130_fd_sc_hd__mux2_1 _10924_ (.A0(_05452_),
    .A1(\data_array.data1[6][16] ),
    .S(_05598_),
    .X(_02669_));
 sky130_fd_sc_hd__mux2_1 _10925_ (.A0(_05454_),
    .A1(\data_array.data1[6][17] ),
    .S(_05598_),
    .X(_02670_));
 sky130_fd_sc_hd__mux2_1 _10926_ (.A0(_05456_),
    .A1(\data_array.data1[6][18] ),
    .S(_05598_),
    .X(_02671_));
 sky130_fd_sc_hd__mux2_1 _10927_ (.A0(_05458_),
    .A1(\data_array.data1[6][19] ),
    .S(_05598_),
    .X(_02672_));
 sky130_fd_sc_hd__mux2_1 _10928_ (.A0(_05460_),
    .A1(\data_array.data1[6][20] ),
    .S(_05598_),
    .X(_02673_));
 sky130_fd_sc_hd__mux2_1 _10929_ (.A0(_05462_),
    .A1(\data_array.data1[6][21] ),
    .S(_05598_),
    .X(_02674_));
 sky130_fd_sc_hd__mux2_1 _10930_ (.A0(_05464_),
    .A1(\data_array.data1[6][22] ),
    .S(_05598_),
    .X(_02675_));
 sky130_fd_sc_hd__mux2_1 _10931_ (.A0(_05466_),
    .A1(\data_array.data1[6][23] ),
    .S(_05598_),
    .X(_02676_));
 sky130_fd_sc_hd__mux2_1 _10932_ (.A0(_05468_),
    .A1(\data_array.data1[6][24] ),
    .S(_05598_),
    .X(_02677_));
 sky130_fd_sc_hd__mux2_1 _10933_ (.A0(_05470_),
    .A1(\data_array.data1[6][25] ),
    .S(_05598_),
    .X(_02678_));
 sky130_fd_sc_hd__mux2_1 _10934_ (.A0(_05472_),
    .A1(\data_array.data1[6][26] ),
    .S(_05598_),
    .X(_02679_));
 sky130_fd_sc_hd__mux2_1 _10935_ (.A0(_05474_),
    .A1(\data_array.data1[6][27] ),
    .S(_05598_),
    .X(_02680_));
 sky130_fd_sc_hd__mux2_1 _10936_ (.A0(_05476_),
    .A1(\data_array.data1[6][28] ),
    .S(_05598_),
    .X(_02681_));
 sky130_fd_sc_hd__mux2_1 _10937_ (.A0(_05478_),
    .A1(\data_array.data1[6][29] ),
    .S(_05598_),
    .X(_02682_));
 sky130_fd_sc_hd__mux2_1 _10938_ (.A0(_05480_),
    .A1(\data_array.data1[6][30] ),
    .S(_05598_),
    .X(_02683_));
 sky130_fd_sc_hd__mux2_1 _10939_ (.A0(_05482_),
    .A1(\data_array.data1[6][31] ),
    .S(_05598_),
    .X(_02684_));
 sky130_fd_sc_hd__mux2_1 _10940_ (.A0(_05484_),
    .A1(\data_array.data1[6][32] ),
    .S(_05598_),
    .X(_02685_));
 sky130_fd_sc_hd__mux2_1 _10941_ (.A0(_05486_),
    .A1(\data_array.data1[6][33] ),
    .S(_05598_),
    .X(_02686_));
 sky130_fd_sc_hd__mux2_1 _10942_ (.A0(_05488_),
    .A1(\data_array.data1[6][34] ),
    .S(_05598_),
    .X(_02687_));
 sky130_fd_sc_hd__mux2_1 _10943_ (.A0(_05490_),
    .A1(\data_array.data1[6][35] ),
    .S(_05598_),
    .X(_02688_));
 sky130_fd_sc_hd__mux2_1 _10944_ (.A0(_05492_),
    .A1(\data_array.data1[6][36] ),
    .S(_05598_),
    .X(_02689_));
 sky130_fd_sc_hd__mux2_1 _10945_ (.A0(_05494_),
    .A1(\data_array.data1[6][37] ),
    .S(_05598_),
    .X(_02690_));
 sky130_fd_sc_hd__mux2_1 _10946_ (.A0(_05496_),
    .A1(\data_array.data1[6][38] ),
    .S(_05598_),
    .X(_02691_));
 sky130_fd_sc_hd__mux2_1 _10947_ (.A0(_05498_),
    .A1(\data_array.data1[6][39] ),
    .S(_05598_),
    .X(_02692_));
 sky130_fd_sc_hd__mux2_1 _10948_ (.A0(_05500_),
    .A1(\data_array.data1[6][40] ),
    .S(_05598_),
    .X(_02693_));
 sky130_fd_sc_hd__mux2_1 _10949_ (.A0(_05502_),
    .A1(\data_array.data1[6][41] ),
    .S(_05598_),
    .X(_02694_));
 sky130_fd_sc_hd__mux2_1 _10950_ (.A0(_05504_),
    .A1(\data_array.data1[6][42] ),
    .S(_05598_),
    .X(_02695_));
 sky130_fd_sc_hd__mux2_1 _10951_ (.A0(_05506_),
    .A1(\data_array.data1[6][43] ),
    .S(_05598_),
    .X(_02696_));
 sky130_fd_sc_hd__mux2_1 _10952_ (.A0(_05508_),
    .A1(\data_array.data1[6][44] ),
    .S(_05598_),
    .X(_02697_));
 sky130_fd_sc_hd__mux2_1 _10953_ (.A0(_05510_),
    .A1(\data_array.data1[6][45] ),
    .S(_05598_),
    .X(_02698_));
 sky130_fd_sc_hd__mux2_1 _10954_ (.A0(_05512_),
    .A1(\data_array.data1[6][46] ),
    .S(_05598_),
    .X(_02699_));
 sky130_fd_sc_hd__mux2_1 _10955_ (.A0(_05514_),
    .A1(\data_array.data1[6][47] ),
    .S(_05598_),
    .X(_02700_));
 sky130_fd_sc_hd__mux2_1 _10956_ (.A0(_05516_),
    .A1(\data_array.data1[6][48] ),
    .S(_05598_),
    .X(_02701_));
 sky130_fd_sc_hd__mux2_1 _10957_ (.A0(_05518_),
    .A1(\data_array.data1[6][49] ),
    .S(_05598_),
    .X(_02702_));
 sky130_fd_sc_hd__mux2_1 _10958_ (.A0(_05520_),
    .A1(\data_array.data1[6][50] ),
    .S(_05598_),
    .X(_02703_));
 sky130_fd_sc_hd__mux2_1 _10959_ (.A0(_05522_),
    .A1(\data_array.data1[6][51] ),
    .S(_05598_),
    .X(_02704_));
 sky130_fd_sc_hd__mux2_1 _10960_ (.A0(_05524_),
    .A1(\data_array.data1[6][52] ),
    .S(_05598_),
    .X(_02705_));
 sky130_fd_sc_hd__mux2_1 _10961_ (.A0(_05526_),
    .A1(\data_array.data1[6][53] ),
    .S(_05598_),
    .X(_02706_));
 sky130_fd_sc_hd__mux2_1 _10962_ (.A0(_05528_),
    .A1(\data_array.data1[6][54] ),
    .S(_05598_),
    .X(_02707_));
 sky130_fd_sc_hd__mux2_1 _10963_ (.A0(_05530_),
    .A1(\data_array.data1[6][55] ),
    .S(_05598_),
    .X(_02708_));
 sky130_fd_sc_hd__mux2_1 _10964_ (.A0(_05532_),
    .A1(\data_array.data1[6][56] ),
    .S(_05598_),
    .X(_02709_));
 sky130_fd_sc_hd__mux2_1 _10965_ (.A0(_05534_),
    .A1(\data_array.data1[6][57] ),
    .S(_05598_),
    .X(_02710_));
 sky130_fd_sc_hd__mux2_1 _10966_ (.A0(_05536_),
    .A1(\data_array.data1[6][58] ),
    .S(_05598_),
    .X(_02711_));
 sky130_fd_sc_hd__mux2_1 _10967_ (.A0(_05538_),
    .A1(\data_array.data1[6][59] ),
    .S(_05598_),
    .X(_02712_));
 sky130_fd_sc_hd__mux2_1 _10968_ (.A0(_05540_),
    .A1(\data_array.data1[6][60] ),
    .S(_05598_),
    .X(_02713_));
 sky130_fd_sc_hd__mux2_1 _10969_ (.A0(_05542_),
    .A1(\data_array.data1[6][61] ),
    .S(_05598_),
    .X(_02714_));
 sky130_fd_sc_hd__mux2_1 _10970_ (.A0(_05544_),
    .A1(\data_array.data1[6][62] ),
    .S(_05598_),
    .X(_02715_));
 sky130_fd_sc_hd__mux2_1 _10971_ (.A0(_05546_),
    .A1(\data_array.data1[6][63] ),
    .S(_05598_),
    .X(_02716_));
 sky130_fd_sc_hd__and2_2 _10972_ (.A(_05415_),
    .B(_05587_),
    .X(_03132_));
 sky130_fd_sc_hd__mux2_1 _10973_ (.A0(\data_array.data0[1][0] ),
    .A1(_05420_),
    .S(_03132_),
    .X(_02717_));
 sky130_fd_sc_hd__mux2_1 _10974_ (.A0(\data_array.data0[1][1] ),
    .A1(_05422_),
    .S(_03132_),
    .X(_02718_));
 sky130_fd_sc_hd__mux2_1 _10975_ (.A0(\data_array.data0[1][2] ),
    .A1(_05424_),
    .S(_03132_),
    .X(_02719_));
 sky130_fd_sc_hd__mux2_1 _10976_ (.A0(\data_array.data0[1][3] ),
    .A1(_05426_),
    .S(_03132_),
    .X(_02720_));
 sky130_fd_sc_hd__mux2_1 _10977_ (.A0(\data_array.data0[1][4] ),
    .A1(_05428_),
    .S(_03132_),
    .X(_02721_));
 sky130_fd_sc_hd__mux2_1 _10978_ (.A0(\data_array.data0[1][5] ),
    .A1(_05430_),
    .S(_03132_),
    .X(_02722_));
 sky130_fd_sc_hd__mux2_1 _10979_ (.A0(\data_array.data0[1][6] ),
    .A1(_05432_),
    .S(_03132_),
    .X(_02723_));
 sky130_fd_sc_hd__mux2_1 _10980_ (.A0(\data_array.data0[1][7] ),
    .A1(_05434_),
    .S(_03132_),
    .X(_02724_));
 sky130_fd_sc_hd__mux2_1 _10981_ (.A0(\data_array.data0[1][8] ),
    .A1(_05436_),
    .S(_03132_),
    .X(_02725_));
 sky130_fd_sc_hd__mux2_1 _10982_ (.A0(\data_array.data0[1][9] ),
    .A1(_05438_),
    .S(_03132_),
    .X(_02726_));
 sky130_fd_sc_hd__mux2_1 _10983_ (.A0(\data_array.data0[1][10] ),
    .A1(_05440_),
    .S(_03132_),
    .X(_02727_));
 sky130_fd_sc_hd__mux2_1 _10984_ (.A0(\data_array.data0[1][11] ),
    .A1(_05442_),
    .S(_03132_),
    .X(_02728_));
 sky130_fd_sc_hd__mux2_1 _10985_ (.A0(\data_array.data0[1][12] ),
    .A1(_05444_),
    .S(_03132_),
    .X(_02729_));
 sky130_fd_sc_hd__mux2_1 _10986_ (.A0(\data_array.data0[1][13] ),
    .A1(_05446_),
    .S(_03132_),
    .X(_02730_));
 sky130_fd_sc_hd__mux2_1 _10987_ (.A0(\data_array.data0[1][14] ),
    .A1(_05448_),
    .S(_03132_),
    .X(_02731_));
 sky130_fd_sc_hd__mux2_1 _10988_ (.A0(\data_array.data0[1][15] ),
    .A1(_05450_),
    .S(_03132_),
    .X(_02732_));
 sky130_fd_sc_hd__mux2_1 _10989_ (.A0(\data_array.data0[1][16] ),
    .A1(_05452_),
    .S(_03132_),
    .X(_02733_));
 sky130_fd_sc_hd__mux2_1 _10990_ (.A0(\data_array.data0[1][17] ),
    .A1(_05454_),
    .S(_03132_),
    .X(_02734_));
 sky130_fd_sc_hd__mux2_1 _10991_ (.A0(\data_array.data0[1][18] ),
    .A1(_05456_),
    .S(_03132_),
    .X(_02735_));
 sky130_fd_sc_hd__mux2_1 _10992_ (.A0(\data_array.data0[1][19] ),
    .A1(_05458_),
    .S(_03132_),
    .X(_02736_));
 sky130_fd_sc_hd__mux2_1 _10993_ (.A0(\data_array.data0[1][20] ),
    .A1(_05460_),
    .S(_03132_),
    .X(_02737_));
 sky130_fd_sc_hd__mux2_1 _10994_ (.A0(\data_array.data0[1][21] ),
    .A1(_05462_),
    .S(_03132_),
    .X(_02738_));
 sky130_fd_sc_hd__mux2_1 _10995_ (.A0(\data_array.data0[1][22] ),
    .A1(_05464_),
    .S(_03132_),
    .X(_02739_));
 sky130_fd_sc_hd__mux2_1 _10996_ (.A0(\data_array.data0[1][23] ),
    .A1(_05466_),
    .S(_03132_),
    .X(_02740_));
 sky130_fd_sc_hd__mux2_1 _10997_ (.A0(\data_array.data0[1][24] ),
    .A1(_05468_),
    .S(_03132_),
    .X(_02741_));
 sky130_fd_sc_hd__mux2_1 _10998_ (.A0(\data_array.data0[1][25] ),
    .A1(_05470_),
    .S(_03132_),
    .X(_02742_));
 sky130_fd_sc_hd__mux2_1 _10999_ (.A0(\data_array.data0[1][26] ),
    .A1(_05472_),
    .S(_03132_),
    .X(_02743_));
 sky130_fd_sc_hd__mux2_1 _11000_ (.A0(\data_array.data0[1][27] ),
    .A1(_05474_),
    .S(_03132_),
    .X(_02744_));
 sky130_fd_sc_hd__mux2_1 _11001_ (.A0(\data_array.data0[1][28] ),
    .A1(_05476_),
    .S(_03132_),
    .X(_02745_));
 sky130_fd_sc_hd__mux2_1 _11002_ (.A0(\data_array.data0[1][29] ),
    .A1(_05478_),
    .S(_03132_),
    .X(_02746_));
 sky130_fd_sc_hd__mux2_1 _11003_ (.A0(\data_array.data0[1][30] ),
    .A1(_05480_),
    .S(_03132_),
    .X(_02747_));
 sky130_fd_sc_hd__mux2_1 _11004_ (.A0(\data_array.data0[1][31] ),
    .A1(_05482_),
    .S(_03132_),
    .X(_02748_));
 sky130_fd_sc_hd__mux2_1 _11005_ (.A0(\data_array.data0[1][32] ),
    .A1(_05484_),
    .S(_03132_),
    .X(_02749_));
 sky130_fd_sc_hd__mux2_1 _11006_ (.A0(\data_array.data0[1][33] ),
    .A1(_05486_),
    .S(_03132_),
    .X(_02750_));
 sky130_fd_sc_hd__mux2_1 _11007_ (.A0(\data_array.data0[1][34] ),
    .A1(_05488_),
    .S(_03132_),
    .X(_02751_));
 sky130_fd_sc_hd__mux2_1 _11008_ (.A0(\data_array.data0[1][35] ),
    .A1(_05490_),
    .S(_03132_),
    .X(_02752_));
 sky130_fd_sc_hd__mux2_1 _11009_ (.A0(\data_array.data0[1][36] ),
    .A1(_05492_),
    .S(_03132_),
    .X(_02753_));
 sky130_fd_sc_hd__mux2_1 _11010_ (.A0(\data_array.data0[1][37] ),
    .A1(_05494_),
    .S(_03132_),
    .X(_02754_));
 sky130_fd_sc_hd__mux2_1 _11011_ (.A0(\data_array.data0[1][38] ),
    .A1(_05496_),
    .S(_03132_),
    .X(_02755_));
 sky130_fd_sc_hd__mux2_1 _11012_ (.A0(\data_array.data0[1][39] ),
    .A1(_05498_),
    .S(_03132_),
    .X(_02756_));
 sky130_fd_sc_hd__mux2_1 _11013_ (.A0(\data_array.data0[1][40] ),
    .A1(_05500_),
    .S(_03132_),
    .X(_02757_));
 sky130_fd_sc_hd__mux2_1 _11014_ (.A0(\data_array.data0[1][41] ),
    .A1(_05502_),
    .S(_03132_),
    .X(_02758_));
 sky130_fd_sc_hd__mux2_1 _11015_ (.A0(\data_array.data0[1][42] ),
    .A1(_05504_),
    .S(_03132_),
    .X(_02759_));
 sky130_fd_sc_hd__mux2_1 _11016_ (.A0(\data_array.data0[1][43] ),
    .A1(_05506_),
    .S(_03132_),
    .X(_02760_));
 sky130_fd_sc_hd__mux2_1 _11017_ (.A0(\data_array.data0[1][44] ),
    .A1(_05508_),
    .S(_03132_),
    .X(_02761_));
 sky130_fd_sc_hd__mux2_1 _11018_ (.A0(\data_array.data0[1][45] ),
    .A1(_05510_),
    .S(_03132_),
    .X(_02762_));
 sky130_fd_sc_hd__mux2_1 _11019_ (.A0(\data_array.data0[1][46] ),
    .A1(_05512_),
    .S(_03132_),
    .X(_02763_));
 sky130_fd_sc_hd__mux2_1 _11020_ (.A0(\data_array.data0[1][47] ),
    .A1(_05514_),
    .S(_03132_),
    .X(_02764_));
 sky130_fd_sc_hd__mux2_1 _11021_ (.A0(\data_array.data0[1][48] ),
    .A1(_05516_),
    .S(_03132_),
    .X(_02765_));
 sky130_fd_sc_hd__mux2_1 _11022_ (.A0(\data_array.data0[1][49] ),
    .A1(_05518_),
    .S(_03132_),
    .X(_02766_));
 sky130_fd_sc_hd__mux2_1 _11023_ (.A0(\data_array.data0[1][50] ),
    .A1(_05520_),
    .S(_03132_),
    .X(_02767_));
 sky130_fd_sc_hd__mux2_1 _11024_ (.A0(\data_array.data0[1][51] ),
    .A1(_05522_),
    .S(_03132_),
    .X(_02768_));
 sky130_fd_sc_hd__mux2_1 _11025_ (.A0(\data_array.data0[1][52] ),
    .A1(_05524_),
    .S(_03132_),
    .X(_02769_));
 sky130_fd_sc_hd__mux2_1 _11026_ (.A0(\data_array.data0[1][53] ),
    .A1(_05526_),
    .S(_03132_),
    .X(_02770_));
 sky130_fd_sc_hd__mux2_1 _11027_ (.A0(\data_array.data0[1][54] ),
    .A1(_05528_),
    .S(_03132_),
    .X(_02771_));
 sky130_fd_sc_hd__mux2_1 _11028_ (.A0(\data_array.data0[1][55] ),
    .A1(_05530_),
    .S(_03132_),
    .X(_02772_));
 sky130_fd_sc_hd__mux2_1 _11029_ (.A0(\data_array.data0[1][56] ),
    .A1(_05532_),
    .S(_03132_),
    .X(_02773_));
 sky130_fd_sc_hd__mux2_1 _11030_ (.A0(\data_array.data0[1][57] ),
    .A1(_05534_),
    .S(_03132_),
    .X(_02774_));
 sky130_fd_sc_hd__mux2_1 _11031_ (.A0(\data_array.data0[1][58] ),
    .A1(_05536_),
    .S(_03132_),
    .X(_02775_));
 sky130_fd_sc_hd__mux2_1 _11032_ (.A0(\data_array.data0[1][59] ),
    .A1(_05538_),
    .S(_03132_),
    .X(_02776_));
 sky130_fd_sc_hd__mux2_1 _11033_ (.A0(\data_array.data0[1][60] ),
    .A1(_05540_),
    .S(_03132_),
    .X(_02777_));
 sky130_fd_sc_hd__mux2_1 _11034_ (.A0(\data_array.data0[1][61] ),
    .A1(_05542_),
    .S(_03132_),
    .X(_02778_));
 sky130_fd_sc_hd__mux2_1 _11035_ (.A0(\data_array.data0[1][62] ),
    .A1(_05544_),
    .S(_03132_),
    .X(_02779_));
 sky130_fd_sc_hd__mux2_1 _11036_ (.A0(\data_array.data0[1][63] ),
    .A1(_05546_),
    .S(_03132_),
    .X(_02780_));
 sky130_fd_sc_hd__and2_2 _11037_ (.A(_05352_),
    .B(_05415_),
    .X(_03133_));
 sky130_fd_sc_hd__mux2_1 _11038_ (.A0(\data_array.data0[2][0] ),
    .A1(_05420_),
    .S(_03133_),
    .X(_02781_));
 sky130_fd_sc_hd__mux2_1 _11039_ (.A0(\data_array.data0[2][1] ),
    .A1(_05422_),
    .S(_03133_),
    .X(_02782_));
 sky130_fd_sc_hd__mux2_1 _11040_ (.A0(\data_array.data0[2][2] ),
    .A1(_05424_),
    .S(_03133_),
    .X(_02783_));
 sky130_fd_sc_hd__mux2_1 _11041_ (.A0(\data_array.data0[2][3] ),
    .A1(_05426_),
    .S(_03133_),
    .X(_02784_));
 sky130_fd_sc_hd__mux2_1 _11042_ (.A0(\data_array.data0[2][4] ),
    .A1(_05428_),
    .S(_03133_),
    .X(_02785_));
 sky130_fd_sc_hd__mux2_1 _11043_ (.A0(\data_array.data0[2][5] ),
    .A1(_05430_),
    .S(_03133_),
    .X(_02786_));
 sky130_fd_sc_hd__mux2_1 _11044_ (.A0(\data_array.data0[2][6] ),
    .A1(_05432_),
    .S(_03133_),
    .X(_02787_));
 sky130_fd_sc_hd__mux2_1 _11045_ (.A0(\data_array.data0[2][7] ),
    .A1(_05434_),
    .S(_03133_),
    .X(_02788_));
 sky130_fd_sc_hd__mux2_1 _11046_ (.A0(\data_array.data0[2][8] ),
    .A1(_05436_),
    .S(_03133_),
    .X(_02789_));
 sky130_fd_sc_hd__mux2_1 _11047_ (.A0(\data_array.data0[2][9] ),
    .A1(_05438_),
    .S(_03133_),
    .X(_02790_));
 sky130_fd_sc_hd__mux2_1 _11048_ (.A0(\data_array.data0[2][10] ),
    .A1(_05440_),
    .S(_03133_),
    .X(_02791_));
 sky130_fd_sc_hd__mux2_1 _11049_ (.A0(\data_array.data0[2][11] ),
    .A1(_05442_),
    .S(_03133_),
    .X(_02792_));
 sky130_fd_sc_hd__mux2_1 _11050_ (.A0(\data_array.data0[2][12] ),
    .A1(_05444_),
    .S(_03133_),
    .X(_02793_));
 sky130_fd_sc_hd__mux2_1 _11051_ (.A0(\data_array.data0[2][13] ),
    .A1(_05446_),
    .S(_03133_),
    .X(_02794_));
 sky130_fd_sc_hd__mux2_1 _11052_ (.A0(\data_array.data0[2][14] ),
    .A1(_05448_),
    .S(_03133_),
    .X(_02795_));
 sky130_fd_sc_hd__mux2_1 _11053_ (.A0(\data_array.data0[2][15] ),
    .A1(_05450_),
    .S(_03133_),
    .X(_02796_));
 sky130_fd_sc_hd__mux2_1 _11054_ (.A0(\data_array.data0[2][16] ),
    .A1(_05452_),
    .S(_03133_),
    .X(_02797_));
 sky130_fd_sc_hd__mux2_1 _11055_ (.A0(\data_array.data0[2][17] ),
    .A1(_05454_),
    .S(_03133_),
    .X(_02798_));
 sky130_fd_sc_hd__mux2_1 _11056_ (.A0(\data_array.data0[2][18] ),
    .A1(_05456_),
    .S(_03133_),
    .X(_02799_));
 sky130_fd_sc_hd__mux2_1 _11057_ (.A0(\data_array.data0[2][19] ),
    .A1(_05458_),
    .S(_03133_),
    .X(_02800_));
 sky130_fd_sc_hd__mux2_1 _11058_ (.A0(\data_array.data0[2][20] ),
    .A1(_05460_),
    .S(_03133_),
    .X(_02801_));
 sky130_fd_sc_hd__mux2_1 _11059_ (.A0(\data_array.data0[2][21] ),
    .A1(_05462_),
    .S(_03133_),
    .X(_02802_));
 sky130_fd_sc_hd__mux2_1 _11060_ (.A0(\data_array.data0[2][22] ),
    .A1(_05464_),
    .S(_03133_),
    .X(_02803_));
 sky130_fd_sc_hd__mux2_1 _11061_ (.A0(\data_array.data0[2][23] ),
    .A1(_05466_),
    .S(_03133_),
    .X(_02804_));
 sky130_fd_sc_hd__mux2_1 _11062_ (.A0(\data_array.data0[2][24] ),
    .A1(_05468_),
    .S(_03133_),
    .X(_02805_));
 sky130_fd_sc_hd__mux2_1 _11063_ (.A0(\data_array.data0[2][25] ),
    .A1(_05470_),
    .S(_03133_),
    .X(_02806_));
 sky130_fd_sc_hd__mux2_1 _11064_ (.A0(\data_array.data0[2][26] ),
    .A1(_05472_),
    .S(_03133_),
    .X(_02807_));
 sky130_fd_sc_hd__mux2_1 _11065_ (.A0(\data_array.data0[2][27] ),
    .A1(_05474_),
    .S(_03133_),
    .X(_02808_));
 sky130_fd_sc_hd__mux2_1 _11066_ (.A0(\data_array.data0[2][28] ),
    .A1(_05476_),
    .S(_03133_),
    .X(_02809_));
 sky130_fd_sc_hd__mux2_1 _11067_ (.A0(\data_array.data0[2][29] ),
    .A1(_05478_),
    .S(_03133_),
    .X(_02810_));
 sky130_fd_sc_hd__mux2_1 _11068_ (.A0(\data_array.data0[2][30] ),
    .A1(_05480_),
    .S(_03133_),
    .X(_02811_));
 sky130_fd_sc_hd__mux2_1 _11069_ (.A0(\data_array.data0[2][31] ),
    .A1(_05482_),
    .S(_03133_),
    .X(_02812_));
 sky130_fd_sc_hd__mux2_1 _11070_ (.A0(\data_array.data0[2][32] ),
    .A1(_05484_),
    .S(_03133_),
    .X(_02813_));
 sky130_fd_sc_hd__mux2_1 _11071_ (.A0(\data_array.data0[2][33] ),
    .A1(_05486_),
    .S(_03133_),
    .X(_02814_));
 sky130_fd_sc_hd__mux2_1 _11072_ (.A0(\data_array.data0[2][34] ),
    .A1(_05488_),
    .S(_03133_),
    .X(_02815_));
 sky130_fd_sc_hd__mux2_1 _11073_ (.A0(\data_array.data0[2][35] ),
    .A1(_05490_),
    .S(_03133_),
    .X(_02816_));
 sky130_fd_sc_hd__mux2_1 _11074_ (.A0(\data_array.data0[2][36] ),
    .A1(_05492_),
    .S(_03133_),
    .X(_02817_));
 sky130_fd_sc_hd__mux2_1 _11075_ (.A0(\data_array.data0[2][37] ),
    .A1(_05494_),
    .S(_03133_),
    .X(_02818_));
 sky130_fd_sc_hd__mux2_1 _11076_ (.A0(\data_array.data0[2][38] ),
    .A1(_05496_),
    .S(_03133_),
    .X(_02819_));
 sky130_fd_sc_hd__mux2_1 _11077_ (.A0(\data_array.data0[2][39] ),
    .A1(_05498_),
    .S(_03133_),
    .X(_02820_));
 sky130_fd_sc_hd__mux2_1 _11078_ (.A0(\data_array.data0[2][40] ),
    .A1(_05500_),
    .S(_03133_),
    .X(_02821_));
 sky130_fd_sc_hd__mux2_1 _11079_ (.A0(\data_array.data0[2][41] ),
    .A1(_05502_),
    .S(_03133_),
    .X(_02822_));
 sky130_fd_sc_hd__mux2_1 _11080_ (.A0(\data_array.data0[2][42] ),
    .A1(_05504_),
    .S(_03133_),
    .X(_02823_));
 sky130_fd_sc_hd__mux2_1 _11081_ (.A0(\data_array.data0[2][43] ),
    .A1(_05506_),
    .S(_03133_),
    .X(_02824_));
 sky130_fd_sc_hd__mux2_1 _11082_ (.A0(\data_array.data0[2][44] ),
    .A1(_05508_),
    .S(_03133_),
    .X(_02825_));
 sky130_fd_sc_hd__mux2_1 _11083_ (.A0(\data_array.data0[2][45] ),
    .A1(_05510_),
    .S(_03133_),
    .X(_02826_));
 sky130_fd_sc_hd__mux2_1 _11084_ (.A0(\data_array.data0[2][46] ),
    .A1(_05512_),
    .S(_03133_),
    .X(_02827_));
 sky130_fd_sc_hd__mux2_1 _11085_ (.A0(\data_array.data0[2][47] ),
    .A1(_05514_),
    .S(_03133_),
    .X(_02828_));
 sky130_fd_sc_hd__mux2_1 _11086_ (.A0(\data_array.data0[2][48] ),
    .A1(_05516_),
    .S(_03133_),
    .X(_02829_));
 sky130_fd_sc_hd__mux2_1 _11087_ (.A0(\data_array.data0[2][49] ),
    .A1(_05518_),
    .S(_03133_),
    .X(_02830_));
 sky130_fd_sc_hd__mux2_1 _11088_ (.A0(\data_array.data0[2][50] ),
    .A1(_05520_),
    .S(_03133_),
    .X(_02831_));
 sky130_fd_sc_hd__mux2_1 _11089_ (.A0(\data_array.data0[2][51] ),
    .A1(_05522_),
    .S(_03133_),
    .X(_02832_));
 sky130_fd_sc_hd__mux2_1 _11090_ (.A0(\data_array.data0[2][52] ),
    .A1(_05524_),
    .S(_03133_),
    .X(_02833_));
 sky130_fd_sc_hd__mux2_1 _11091_ (.A0(\data_array.data0[2][53] ),
    .A1(_05526_),
    .S(_03133_),
    .X(_02834_));
 sky130_fd_sc_hd__mux2_1 _11092_ (.A0(\data_array.data0[2][54] ),
    .A1(_05528_),
    .S(_03133_),
    .X(_02835_));
 sky130_fd_sc_hd__mux2_1 _11093_ (.A0(\data_array.data0[2][55] ),
    .A1(_05530_),
    .S(_03133_),
    .X(_02836_));
 sky130_fd_sc_hd__mux2_1 _11094_ (.A0(\data_array.data0[2][56] ),
    .A1(_05532_),
    .S(_03133_),
    .X(_02837_));
 sky130_fd_sc_hd__mux2_1 _11095_ (.A0(\data_array.data0[2][57] ),
    .A1(_05534_),
    .S(_03133_),
    .X(_02838_));
 sky130_fd_sc_hd__mux2_1 _11096_ (.A0(\data_array.data0[2][58] ),
    .A1(_05536_),
    .S(_03133_),
    .X(_02839_));
 sky130_fd_sc_hd__mux2_1 _11097_ (.A0(\data_array.data0[2][59] ),
    .A1(_05538_),
    .S(_03133_),
    .X(_02840_));
 sky130_fd_sc_hd__mux2_1 _11098_ (.A0(\data_array.data0[2][60] ),
    .A1(_05540_),
    .S(_03133_),
    .X(_02841_));
 sky130_fd_sc_hd__mux2_1 _11099_ (.A0(\data_array.data0[2][61] ),
    .A1(_05542_),
    .S(_03133_),
    .X(_02842_));
 sky130_fd_sc_hd__mux2_1 _11100_ (.A0(\data_array.data0[2][62] ),
    .A1(_05544_),
    .S(_03133_),
    .X(_02843_));
 sky130_fd_sc_hd__mux2_1 _11101_ (.A0(\data_array.data0[2][63] ),
    .A1(_05546_),
    .S(_03133_),
    .X(_02844_));
 sky130_fd_sc_hd__mux2_1 _11102_ (.A0(_05420_),
    .A1(\data_array.data1[12][0] ),
    .S(_05594_),
    .X(_02845_));
 sky130_fd_sc_hd__mux2_1 _11103_ (.A0(_05422_),
    .A1(\data_array.data1[12][1] ),
    .S(_05594_),
    .X(_02846_));
 sky130_fd_sc_hd__mux2_1 _11104_ (.A0(_05424_),
    .A1(\data_array.data1[12][2] ),
    .S(_05594_),
    .X(_02847_));
 sky130_fd_sc_hd__mux2_1 _11105_ (.A0(_05426_),
    .A1(\data_array.data1[12][3] ),
    .S(_05594_),
    .X(_02848_));
 sky130_fd_sc_hd__mux2_1 _11106_ (.A0(_05428_),
    .A1(\data_array.data1[12][4] ),
    .S(_05594_),
    .X(_02849_));
 sky130_fd_sc_hd__mux2_1 _11107_ (.A0(_05430_),
    .A1(\data_array.data1[12][5] ),
    .S(_05594_),
    .X(_02850_));
 sky130_fd_sc_hd__mux2_1 _11108_ (.A0(_05432_),
    .A1(\data_array.data1[12][6] ),
    .S(_05594_),
    .X(_02851_));
 sky130_fd_sc_hd__mux2_1 _11109_ (.A0(_05434_),
    .A1(\data_array.data1[12][7] ),
    .S(_05594_),
    .X(_02852_));
 sky130_fd_sc_hd__mux2_1 _11110_ (.A0(_05436_),
    .A1(\data_array.data1[12][8] ),
    .S(_05594_),
    .X(_02853_));
 sky130_fd_sc_hd__mux2_1 _11111_ (.A0(_05438_),
    .A1(\data_array.data1[12][9] ),
    .S(_05594_),
    .X(_02854_));
 sky130_fd_sc_hd__mux2_1 _11112_ (.A0(_05440_),
    .A1(\data_array.data1[12][10] ),
    .S(_05594_),
    .X(_02855_));
 sky130_fd_sc_hd__mux2_1 _11113_ (.A0(_05442_),
    .A1(\data_array.data1[12][11] ),
    .S(_05594_),
    .X(_02856_));
 sky130_fd_sc_hd__mux2_1 _11114_ (.A0(_05444_),
    .A1(\data_array.data1[12][12] ),
    .S(_05594_),
    .X(_02857_));
 sky130_fd_sc_hd__mux2_1 _11115_ (.A0(_05446_),
    .A1(\data_array.data1[12][13] ),
    .S(_05594_),
    .X(_02858_));
 sky130_fd_sc_hd__mux2_1 _11116_ (.A0(_05448_),
    .A1(\data_array.data1[12][14] ),
    .S(_05594_),
    .X(_02859_));
 sky130_fd_sc_hd__mux2_1 _11117_ (.A0(_05450_),
    .A1(\data_array.data1[12][15] ),
    .S(_05594_),
    .X(_02860_));
 sky130_fd_sc_hd__mux2_1 _11118_ (.A0(_05452_),
    .A1(\data_array.data1[12][16] ),
    .S(_05594_),
    .X(_02861_));
 sky130_fd_sc_hd__mux2_1 _11119_ (.A0(_05454_),
    .A1(\data_array.data1[12][17] ),
    .S(_05594_),
    .X(_02862_));
 sky130_fd_sc_hd__mux2_1 _11120_ (.A0(_05456_),
    .A1(\data_array.data1[12][18] ),
    .S(_05594_),
    .X(_02863_));
 sky130_fd_sc_hd__mux2_1 _11121_ (.A0(_05458_),
    .A1(\data_array.data1[12][19] ),
    .S(_05594_),
    .X(_02864_));
 sky130_fd_sc_hd__mux2_1 _11122_ (.A0(_05460_),
    .A1(\data_array.data1[12][20] ),
    .S(_05594_),
    .X(_02865_));
 sky130_fd_sc_hd__mux2_1 _11123_ (.A0(_05462_),
    .A1(\data_array.data1[12][21] ),
    .S(_05594_),
    .X(_02866_));
 sky130_fd_sc_hd__mux2_1 _11124_ (.A0(_05464_),
    .A1(\data_array.data1[12][22] ),
    .S(_05594_),
    .X(_02867_));
 sky130_fd_sc_hd__mux2_1 _11125_ (.A0(_05466_),
    .A1(\data_array.data1[12][23] ),
    .S(_05594_),
    .X(_02868_));
 sky130_fd_sc_hd__mux2_1 _11126_ (.A0(_05468_),
    .A1(\data_array.data1[12][24] ),
    .S(_05594_),
    .X(_02869_));
 sky130_fd_sc_hd__mux2_1 _11127_ (.A0(_05470_),
    .A1(\data_array.data1[12][25] ),
    .S(_05594_),
    .X(_02870_));
 sky130_fd_sc_hd__mux2_1 _11128_ (.A0(_05472_),
    .A1(\data_array.data1[12][26] ),
    .S(_05594_),
    .X(_02871_));
 sky130_fd_sc_hd__mux2_1 _11129_ (.A0(_05474_),
    .A1(\data_array.data1[12][27] ),
    .S(_05594_),
    .X(_02872_));
 sky130_fd_sc_hd__mux2_1 _11130_ (.A0(_05476_),
    .A1(\data_array.data1[12][28] ),
    .S(_05594_),
    .X(_02873_));
 sky130_fd_sc_hd__mux2_1 _11131_ (.A0(_05478_),
    .A1(\data_array.data1[12][29] ),
    .S(_05594_),
    .X(_02874_));
 sky130_fd_sc_hd__mux2_1 _11132_ (.A0(_05480_),
    .A1(\data_array.data1[12][30] ),
    .S(_05594_),
    .X(_02875_));
 sky130_fd_sc_hd__mux2_1 _11133_ (.A0(_05482_),
    .A1(\data_array.data1[12][31] ),
    .S(_05594_),
    .X(_02876_));
 sky130_fd_sc_hd__mux2_1 _11134_ (.A0(_05484_),
    .A1(\data_array.data1[12][32] ),
    .S(_05594_),
    .X(_02877_));
 sky130_fd_sc_hd__mux2_1 _11135_ (.A0(_05486_),
    .A1(\data_array.data1[12][33] ),
    .S(_05594_),
    .X(_02878_));
 sky130_fd_sc_hd__mux2_1 _11136_ (.A0(_05488_),
    .A1(\data_array.data1[12][34] ),
    .S(_05594_),
    .X(_02879_));
 sky130_fd_sc_hd__mux2_1 _11137_ (.A0(_05490_),
    .A1(\data_array.data1[12][35] ),
    .S(_05594_),
    .X(_02880_));
 sky130_fd_sc_hd__mux2_1 _11138_ (.A0(_05492_),
    .A1(\data_array.data1[12][36] ),
    .S(_05594_),
    .X(_02881_));
 sky130_fd_sc_hd__mux2_1 _11139_ (.A0(_05494_),
    .A1(\data_array.data1[12][37] ),
    .S(_05594_),
    .X(_02882_));
 sky130_fd_sc_hd__mux2_1 _11140_ (.A0(_05496_),
    .A1(\data_array.data1[12][38] ),
    .S(_05594_),
    .X(_02883_));
 sky130_fd_sc_hd__mux2_1 _11141_ (.A0(_05498_),
    .A1(\data_array.data1[12][39] ),
    .S(_05594_),
    .X(_02884_));
 sky130_fd_sc_hd__mux2_1 _11142_ (.A0(_05500_),
    .A1(\data_array.data1[12][40] ),
    .S(_05594_),
    .X(_02885_));
 sky130_fd_sc_hd__mux2_1 _11143_ (.A0(_05502_),
    .A1(\data_array.data1[12][41] ),
    .S(_05594_),
    .X(_02886_));
 sky130_fd_sc_hd__mux2_1 _11144_ (.A0(_05504_),
    .A1(\data_array.data1[12][42] ),
    .S(_05594_),
    .X(_02887_));
 sky130_fd_sc_hd__mux2_1 _11145_ (.A0(_05506_),
    .A1(\data_array.data1[12][43] ),
    .S(_05594_),
    .X(_02888_));
 sky130_fd_sc_hd__mux2_1 _11146_ (.A0(_05508_),
    .A1(\data_array.data1[12][44] ),
    .S(_05594_),
    .X(_02889_));
 sky130_fd_sc_hd__mux2_1 _11147_ (.A0(_05510_),
    .A1(\data_array.data1[12][45] ),
    .S(_05594_),
    .X(_02890_));
 sky130_fd_sc_hd__mux2_1 _11148_ (.A0(_05512_),
    .A1(\data_array.data1[12][46] ),
    .S(_05594_),
    .X(_02891_));
 sky130_fd_sc_hd__mux2_1 _11149_ (.A0(_05514_),
    .A1(\data_array.data1[12][47] ),
    .S(_05594_),
    .X(_02892_));
 sky130_fd_sc_hd__mux2_1 _11150_ (.A0(_05516_),
    .A1(\data_array.data1[12][48] ),
    .S(_05594_),
    .X(_02893_));
 sky130_fd_sc_hd__mux2_1 _11151_ (.A0(_05518_),
    .A1(\data_array.data1[12][49] ),
    .S(_05594_),
    .X(_02894_));
 sky130_fd_sc_hd__mux2_1 _11152_ (.A0(_05520_),
    .A1(\data_array.data1[12][50] ),
    .S(_05594_),
    .X(_02895_));
 sky130_fd_sc_hd__mux2_1 _11153_ (.A0(_05522_),
    .A1(\data_array.data1[12][51] ),
    .S(_05594_),
    .X(_02896_));
 sky130_fd_sc_hd__mux2_1 _11154_ (.A0(_05524_),
    .A1(\data_array.data1[12][52] ),
    .S(_05594_),
    .X(_02897_));
 sky130_fd_sc_hd__mux2_1 _11155_ (.A0(_05526_),
    .A1(\data_array.data1[12][53] ),
    .S(_05594_),
    .X(_02898_));
 sky130_fd_sc_hd__mux2_1 _11156_ (.A0(_05528_),
    .A1(\data_array.data1[12][54] ),
    .S(_05594_),
    .X(_02899_));
 sky130_fd_sc_hd__mux2_1 _11157_ (.A0(_05530_),
    .A1(\data_array.data1[12][55] ),
    .S(_05594_),
    .X(_02900_));
 sky130_fd_sc_hd__mux2_1 _11158_ (.A0(_05532_),
    .A1(\data_array.data1[12][56] ),
    .S(_05594_),
    .X(_02901_));
 sky130_fd_sc_hd__mux2_1 _11159_ (.A0(_05534_),
    .A1(\data_array.data1[12][57] ),
    .S(_05594_),
    .X(_02902_));
 sky130_fd_sc_hd__mux2_1 _11160_ (.A0(_05536_),
    .A1(\data_array.data1[12][58] ),
    .S(_05594_),
    .X(_02903_));
 sky130_fd_sc_hd__mux2_1 _11161_ (.A0(_05538_),
    .A1(\data_array.data1[12][59] ),
    .S(_05594_),
    .X(_02904_));
 sky130_fd_sc_hd__mux2_1 _11162_ (.A0(_05540_),
    .A1(\data_array.data1[12][60] ),
    .S(_05594_),
    .X(_02905_));
 sky130_fd_sc_hd__mux2_1 _11163_ (.A0(_05542_),
    .A1(\data_array.data1[12][61] ),
    .S(_05594_),
    .X(_02906_));
 sky130_fd_sc_hd__mux2_1 _11164_ (.A0(_05544_),
    .A1(\data_array.data1[12][62] ),
    .S(_05594_),
    .X(_02907_));
 sky130_fd_sc_hd__mux2_1 _11165_ (.A0(_05546_),
    .A1(\data_array.data1[12][63] ),
    .S(_05594_),
    .X(_02908_));
 sky130_fd_sc_hd__mux2_1 _11166_ (.A0(_05420_),
    .A1(\data_array.data1[11][0] ),
    .S(_05551_),
    .X(_02909_));
 sky130_fd_sc_hd__mux2_1 _11167_ (.A0(_05422_),
    .A1(\data_array.data1[11][1] ),
    .S(_05551_),
    .X(_02910_));
 sky130_fd_sc_hd__mux2_1 _11168_ (.A0(_05424_),
    .A1(\data_array.data1[11][2] ),
    .S(_05551_),
    .X(_02911_));
 sky130_fd_sc_hd__mux2_1 _11169_ (.A0(_05426_),
    .A1(\data_array.data1[11][3] ),
    .S(_05551_),
    .X(_02912_));
 sky130_fd_sc_hd__mux2_1 _11170_ (.A0(_05428_),
    .A1(\data_array.data1[11][4] ),
    .S(_05551_),
    .X(_02913_));
 sky130_fd_sc_hd__mux2_1 _11171_ (.A0(_05430_),
    .A1(\data_array.data1[11][5] ),
    .S(_05551_),
    .X(_02914_));
 sky130_fd_sc_hd__mux2_1 _11172_ (.A0(_05432_),
    .A1(\data_array.data1[11][6] ),
    .S(_05551_),
    .X(_02915_));
 sky130_fd_sc_hd__mux2_1 _11173_ (.A0(_05434_),
    .A1(\data_array.data1[11][7] ),
    .S(_05551_),
    .X(_02916_));
 sky130_fd_sc_hd__mux2_1 _11174_ (.A0(_05436_),
    .A1(\data_array.data1[11][8] ),
    .S(_05551_),
    .X(_02917_));
 sky130_fd_sc_hd__mux2_1 _11175_ (.A0(_05438_),
    .A1(\data_array.data1[11][9] ),
    .S(_05551_),
    .X(_02918_));
 sky130_fd_sc_hd__mux2_1 _11176_ (.A0(_05440_),
    .A1(\data_array.data1[11][10] ),
    .S(_05551_),
    .X(_02919_));
 sky130_fd_sc_hd__mux2_1 _11177_ (.A0(_05442_),
    .A1(\data_array.data1[11][11] ),
    .S(_05551_),
    .X(_02920_));
 sky130_fd_sc_hd__mux2_1 _11178_ (.A0(_05444_),
    .A1(\data_array.data1[11][12] ),
    .S(_05551_),
    .X(_02921_));
 sky130_fd_sc_hd__mux2_1 _11179_ (.A0(_05446_),
    .A1(\data_array.data1[11][13] ),
    .S(_05551_),
    .X(_02922_));
 sky130_fd_sc_hd__mux2_1 _11180_ (.A0(_05448_),
    .A1(\data_array.data1[11][14] ),
    .S(_05551_),
    .X(_02923_));
 sky130_fd_sc_hd__mux2_1 _11181_ (.A0(_05450_),
    .A1(\data_array.data1[11][15] ),
    .S(_05551_),
    .X(_02924_));
 sky130_fd_sc_hd__mux2_1 _11182_ (.A0(_05452_),
    .A1(\data_array.data1[11][16] ),
    .S(_05551_),
    .X(_02925_));
 sky130_fd_sc_hd__mux2_1 _11183_ (.A0(_05454_),
    .A1(\data_array.data1[11][17] ),
    .S(_05551_),
    .X(_02926_));
 sky130_fd_sc_hd__mux2_1 _11184_ (.A0(_05456_),
    .A1(\data_array.data1[11][18] ),
    .S(_05551_),
    .X(_02927_));
 sky130_fd_sc_hd__mux2_1 _11185_ (.A0(_05458_),
    .A1(\data_array.data1[11][19] ),
    .S(_05551_),
    .X(_02928_));
 sky130_fd_sc_hd__mux2_1 _11186_ (.A0(_05460_),
    .A1(\data_array.data1[11][20] ),
    .S(_05551_),
    .X(_02929_));
 sky130_fd_sc_hd__mux2_1 _11187_ (.A0(_05462_),
    .A1(\data_array.data1[11][21] ),
    .S(_05551_),
    .X(_02930_));
 sky130_fd_sc_hd__mux2_1 _11188_ (.A0(_05464_),
    .A1(\data_array.data1[11][22] ),
    .S(_05551_),
    .X(_02931_));
 sky130_fd_sc_hd__mux2_1 _11189_ (.A0(_05466_),
    .A1(\data_array.data1[11][23] ),
    .S(_05551_),
    .X(_02932_));
 sky130_fd_sc_hd__mux2_1 _11190_ (.A0(_05468_),
    .A1(\data_array.data1[11][24] ),
    .S(_05551_),
    .X(_02933_));
 sky130_fd_sc_hd__mux2_1 _11191_ (.A0(_05470_),
    .A1(\data_array.data1[11][25] ),
    .S(_05551_),
    .X(_02934_));
 sky130_fd_sc_hd__mux2_1 _11192_ (.A0(_05472_),
    .A1(\data_array.data1[11][26] ),
    .S(_05551_),
    .X(_02935_));
 sky130_fd_sc_hd__mux2_1 _11193_ (.A0(_05474_),
    .A1(\data_array.data1[11][27] ),
    .S(_05551_),
    .X(_02936_));
 sky130_fd_sc_hd__mux2_1 _11194_ (.A0(_05476_),
    .A1(\data_array.data1[11][28] ),
    .S(_05551_),
    .X(_02937_));
 sky130_fd_sc_hd__mux2_1 _11195_ (.A0(_05478_),
    .A1(\data_array.data1[11][29] ),
    .S(_05551_),
    .X(_02938_));
 sky130_fd_sc_hd__mux2_1 _11196_ (.A0(_05480_),
    .A1(\data_array.data1[11][30] ),
    .S(_05551_),
    .X(_02939_));
 sky130_fd_sc_hd__mux2_1 _11197_ (.A0(_05482_),
    .A1(\data_array.data1[11][31] ),
    .S(_05551_),
    .X(_02940_));
 sky130_fd_sc_hd__mux2_1 _11198_ (.A0(_05484_),
    .A1(\data_array.data1[11][32] ),
    .S(_05551_),
    .X(_02941_));
 sky130_fd_sc_hd__mux2_1 _11199_ (.A0(_05486_),
    .A1(\data_array.data1[11][33] ),
    .S(_05551_),
    .X(_02942_));
 sky130_fd_sc_hd__mux2_1 _11200_ (.A0(_05488_),
    .A1(\data_array.data1[11][34] ),
    .S(_05551_),
    .X(_02943_));
 sky130_fd_sc_hd__mux2_1 _11201_ (.A0(_05490_),
    .A1(\data_array.data1[11][35] ),
    .S(_05551_),
    .X(_02944_));
 sky130_fd_sc_hd__mux2_1 _11202_ (.A0(_05492_),
    .A1(\data_array.data1[11][36] ),
    .S(_05551_),
    .X(_02945_));
 sky130_fd_sc_hd__mux2_1 _11203_ (.A0(_05494_),
    .A1(\data_array.data1[11][37] ),
    .S(_05551_),
    .X(_02946_));
 sky130_fd_sc_hd__mux2_1 _11204_ (.A0(_05496_),
    .A1(\data_array.data1[11][38] ),
    .S(_05551_),
    .X(_02947_));
 sky130_fd_sc_hd__mux2_1 _11205_ (.A0(_05498_),
    .A1(\data_array.data1[11][39] ),
    .S(_05551_),
    .X(_02948_));
 sky130_fd_sc_hd__mux2_1 _11206_ (.A0(_05500_),
    .A1(\data_array.data1[11][40] ),
    .S(_05551_),
    .X(_02949_));
 sky130_fd_sc_hd__mux2_1 _11207_ (.A0(_05502_),
    .A1(\data_array.data1[11][41] ),
    .S(_05551_),
    .X(_02950_));
 sky130_fd_sc_hd__mux2_1 _11208_ (.A0(_05504_),
    .A1(\data_array.data1[11][42] ),
    .S(_05551_),
    .X(_02951_));
 sky130_fd_sc_hd__mux2_1 _11209_ (.A0(_05506_),
    .A1(\data_array.data1[11][43] ),
    .S(_05551_),
    .X(_02952_));
 sky130_fd_sc_hd__mux2_1 _11210_ (.A0(_05508_),
    .A1(\data_array.data1[11][44] ),
    .S(_05551_),
    .X(_02953_));
 sky130_fd_sc_hd__mux2_1 _11211_ (.A0(_05510_),
    .A1(\data_array.data1[11][45] ),
    .S(_05551_),
    .X(_02954_));
 sky130_fd_sc_hd__mux2_1 _11212_ (.A0(_05512_),
    .A1(\data_array.data1[11][46] ),
    .S(_05551_),
    .X(_02955_));
 sky130_fd_sc_hd__mux2_1 _11213_ (.A0(_05514_),
    .A1(\data_array.data1[11][47] ),
    .S(_05551_),
    .X(_02956_));
 sky130_fd_sc_hd__mux2_1 _11214_ (.A0(_05516_),
    .A1(\data_array.data1[11][48] ),
    .S(_05551_),
    .X(_02957_));
 sky130_fd_sc_hd__mux2_1 _11215_ (.A0(_05518_),
    .A1(\data_array.data1[11][49] ),
    .S(_05551_),
    .X(_02958_));
 sky130_fd_sc_hd__mux2_1 _11216_ (.A0(_05520_),
    .A1(\data_array.data1[11][50] ),
    .S(_05551_),
    .X(_02959_));
 sky130_fd_sc_hd__mux2_1 _11217_ (.A0(_05522_),
    .A1(\data_array.data1[11][51] ),
    .S(_05551_),
    .X(_02960_));
 sky130_fd_sc_hd__mux2_1 _11218_ (.A0(_05524_),
    .A1(\data_array.data1[11][52] ),
    .S(_05551_),
    .X(_02961_));
 sky130_fd_sc_hd__mux2_1 _11219_ (.A0(_05526_),
    .A1(\data_array.data1[11][53] ),
    .S(_05551_),
    .X(_02962_));
 sky130_fd_sc_hd__mux2_1 _11220_ (.A0(_05528_),
    .A1(\data_array.data1[11][54] ),
    .S(_05551_),
    .X(_02963_));
 sky130_fd_sc_hd__mux2_1 _11221_ (.A0(_05530_),
    .A1(\data_array.data1[11][55] ),
    .S(_05551_),
    .X(_02964_));
 sky130_fd_sc_hd__mux2_1 _11222_ (.A0(_05532_),
    .A1(\data_array.data1[11][56] ),
    .S(_05551_),
    .X(_02965_));
 sky130_fd_sc_hd__mux2_1 _11223_ (.A0(_05534_),
    .A1(\data_array.data1[11][57] ),
    .S(_05551_),
    .X(_02966_));
 sky130_fd_sc_hd__mux2_1 _11224_ (.A0(_05536_),
    .A1(\data_array.data1[11][58] ),
    .S(_05551_),
    .X(_02967_));
 sky130_fd_sc_hd__mux2_1 _11225_ (.A0(_05538_),
    .A1(\data_array.data1[11][59] ),
    .S(_05551_),
    .X(_02968_));
 sky130_fd_sc_hd__mux2_1 _11226_ (.A0(_05540_),
    .A1(\data_array.data1[11][60] ),
    .S(_05551_),
    .X(_02969_));
 sky130_fd_sc_hd__mux2_1 _11227_ (.A0(_05542_),
    .A1(\data_array.data1[11][61] ),
    .S(_05551_),
    .X(_02970_));
 sky130_fd_sc_hd__mux2_1 _11228_ (.A0(_05544_),
    .A1(\data_array.data1[11][62] ),
    .S(_05551_),
    .X(_02971_));
 sky130_fd_sc_hd__mux2_1 _11229_ (.A0(_05546_),
    .A1(\data_array.data1[11][63] ),
    .S(_05551_),
    .X(_02972_));
 sky130_fd_sc_hd__mux2_1 _11230_ (.A0(_05420_),
    .A1(\data_array.data1[10][0] ),
    .S(_05548_),
    .X(_02973_));
 sky130_fd_sc_hd__mux2_1 _11231_ (.A0(_05422_),
    .A1(\data_array.data1[10][1] ),
    .S(_05548_),
    .X(_02974_));
 sky130_fd_sc_hd__mux2_1 _11232_ (.A0(_05424_),
    .A1(\data_array.data1[10][2] ),
    .S(_05548_),
    .X(_02975_));
 sky130_fd_sc_hd__mux2_1 _11233_ (.A0(_05426_),
    .A1(\data_array.data1[10][3] ),
    .S(_05548_),
    .X(_02976_));
 sky130_fd_sc_hd__mux2_1 _11234_ (.A0(_05428_),
    .A1(\data_array.data1[10][4] ),
    .S(_05548_),
    .X(_02977_));
 sky130_fd_sc_hd__mux2_1 _11235_ (.A0(_05430_),
    .A1(\data_array.data1[10][5] ),
    .S(_05548_),
    .X(_02978_));
 sky130_fd_sc_hd__mux2_1 _11236_ (.A0(_05432_),
    .A1(\data_array.data1[10][6] ),
    .S(_05548_),
    .X(_02979_));
 sky130_fd_sc_hd__mux2_1 _11237_ (.A0(_05434_),
    .A1(\data_array.data1[10][7] ),
    .S(_05548_),
    .X(_02980_));
 sky130_fd_sc_hd__mux2_1 _11238_ (.A0(_05436_),
    .A1(\data_array.data1[10][8] ),
    .S(_05548_),
    .X(_02981_));
 sky130_fd_sc_hd__mux2_1 _11239_ (.A0(_05438_),
    .A1(\data_array.data1[10][9] ),
    .S(_05548_),
    .X(_02982_));
 sky130_fd_sc_hd__mux2_1 _11240_ (.A0(_05440_),
    .A1(\data_array.data1[10][10] ),
    .S(_05548_),
    .X(_02983_));
 sky130_fd_sc_hd__mux2_1 _11241_ (.A0(_05442_),
    .A1(\data_array.data1[10][11] ),
    .S(_05548_),
    .X(_02984_));
 sky130_fd_sc_hd__mux2_1 _11242_ (.A0(_05444_),
    .A1(\data_array.data1[10][12] ),
    .S(_05548_),
    .X(_02985_));
 sky130_fd_sc_hd__mux2_1 _11243_ (.A0(_05446_),
    .A1(\data_array.data1[10][13] ),
    .S(_05548_),
    .X(_02986_));
 sky130_fd_sc_hd__mux2_1 _11244_ (.A0(_05448_),
    .A1(\data_array.data1[10][14] ),
    .S(_05548_),
    .X(_02987_));
 sky130_fd_sc_hd__mux2_1 _11245_ (.A0(_05450_),
    .A1(\data_array.data1[10][15] ),
    .S(_05548_),
    .X(_02988_));
 sky130_fd_sc_hd__mux2_1 _11246_ (.A0(_05452_),
    .A1(\data_array.data1[10][16] ),
    .S(_05548_),
    .X(_02989_));
 sky130_fd_sc_hd__mux2_1 _11247_ (.A0(_05454_),
    .A1(\data_array.data1[10][17] ),
    .S(_05548_),
    .X(_02990_));
 sky130_fd_sc_hd__mux2_1 _11248_ (.A0(_05456_),
    .A1(\data_array.data1[10][18] ),
    .S(_05548_),
    .X(_02991_));
 sky130_fd_sc_hd__mux2_1 _11249_ (.A0(_05458_),
    .A1(\data_array.data1[10][19] ),
    .S(_05548_),
    .X(_02992_));
 sky130_fd_sc_hd__mux2_1 _11250_ (.A0(_05460_),
    .A1(\data_array.data1[10][20] ),
    .S(_05548_),
    .X(_02993_));
 sky130_fd_sc_hd__mux2_1 _11251_ (.A0(_05462_),
    .A1(\data_array.data1[10][21] ),
    .S(_05548_),
    .X(_02994_));
 sky130_fd_sc_hd__mux2_1 _11252_ (.A0(_05464_),
    .A1(\data_array.data1[10][22] ),
    .S(_05548_),
    .X(_02995_));
 sky130_fd_sc_hd__mux2_1 _11253_ (.A0(_05466_),
    .A1(\data_array.data1[10][23] ),
    .S(_05548_),
    .X(_02996_));
 sky130_fd_sc_hd__mux2_1 _11254_ (.A0(_05468_),
    .A1(\data_array.data1[10][24] ),
    .S(_05548_),
    .X(_02997_));
 sky130_fd_sc_hd__mux2_1 _11255_ (.A0(_05470_),
    .A1(\data_array.data1[10][25] ),
    .S(_05548_),
    .X(_02998_));
 sky130_fd_sc_hd__mux2_1 _11256_ (.A0(_05472_),
    .A1(\data_array.data1[10][26] ),
    .S(_05548_),
    .X(_02999_));
 sky130_fd_sc_hd__mux2_1 _11257_ (.A0(_05474_),
    .A1(\data_array.data1[10][27] ),
    .S(_05548_),
    .X(_03000_));
 sky130_fd_sc_hd__mux2_1 _11258_ (.A0(_05476_),
    .A1(\data_array.data1[10][28] ),
    .S(_05548_),
    .X(_03001_));
 sky130_fd_sc_hd__mux2_1 _11259_ (.A0(_05478_),
    .A1(\data_array.data1[10][29] ),
    .S(_05548_),
    .X(_03002_));
 sky130_fd_sc_hd__mux2_1 _11260_ (.A0(_05480_),
    .A1(\data_array.data1[10][30] ),
    .S(_05548_),
    .X(_03003_));
 sky130_fd_sc_hd__mux2_1 _11261_ (.A0(_05482_),
    .A1(\data_array.data1[10][31] ),
    .S(_05548_),
    .X(_03004_));
 sky130_fd_sc_hd__mux2_1 _11262_ (.A0(_05484_),
    .A1(\data_array.data1[10][32] ),
    .S(_05548_),
    .X(_03005_));
 sky130_fd_sc_hd__mux2_1 _11263_ (.A0(_05486_),
    .A1(\data_array.data1[10][33] ),
    .S(_05548_),
    .X(_03006_));
 sky130_fd_sc_hd__mux2_1 _11264_ (.A0(_05488_),
    .A1(\data_array.data1[10][34] ),
    .S(_05548_),
    .X(_03007_));
 sky130_fd_sc_hd__mux2_1 _11265_ (.A0(_05490_),
    .A1(\data_array.data1[10][35] ),
    .S(_05548_),
    .X(_03008_));
 sky130_fd_sc_hd__mux2_1 _11266_ (.A0(_05492_),
    .A1(\data_array.data1[10][36] ),
    .S(_05548_),
    .X(_03009_));
 sky130_fd_sc_hd__mux2_1 _11267_ (.A0(_05494_),
    .A1(\data_array.data1[10][37] ),
    .S(_05548_),
    .X(_03010_));
 sky130_fd_sc_hd__mux2_1 _11268_ (.A0(_05496_),
    .A1(\data_array.data1[10][38] ),
    .S(_05548_),
    .X(_03011_));
 sky130_fd_sc_hd__mux2_1 _11269_ (.A0(_05498_),
    .A1(\data_array.data1[10][39] ),
    .S(_05548_),
    .X(_03012_));
 sky130_fd_sc_hd__mux2_1 _11270_ (.A0(_05500_),
    .A1(\data_array.data1[10][40] ),
    .S(_05548_),
    .X(_03013_));
 sky130_fd_sc_hd__mux2_1 _11271_ (.A0(_05502_),
    .A1(\data_array.data1[10][41] ),
    .S(_05548_),
    .X(_03014_));
 sky130_fd_sc_hd__mux2_1 _11272_ (.A0(_05504_),
    .A1(\data_array.data1[10][42] ),
    .S(_05548_),
    .X(_03015_));
 sky130_fd_sc_hd__mux2_1 _11273_ (.A0(_05506_),
    .A1(\data_array.data1[10][43] ),
    .S(_05548_),
    .X(_03016_));
 sky130_fd_sc_hd__mux2_1 _11274_ (.A0(_05508_),
    .A1(\data_array.data1[10][44] ),
    .S(_05548_),
    .X(_03017_));
 sky130_fd_sc_hd__mux2_1 _11275_ (.A0(_05510_),
    .A1(\data_array.data1[10][45] ),
    .S(_05548_),
    .X(_03018_));
 sky130_fd_sc_hd__mux2_1 _11276_ (.A0(_05512_),
    .A1(\data_array.data1[10][46] ),
    .S(_05548_),
    .X(_03019_));
 sky130_fd_sc_hd__mux2_1 _11277_ (.A0(_05514_),
    .A1(\data_array.data1[10][47] ),
    .S(_05548_),
    .X(_03020_));
 sky130_fd_sc_hd__mux2_1 _11278_ (.A0(_05516_),
    .A1(\data_array.data1[10][48] ),
    .S(_05548_),
    .X(_03021_));
 sky130_fd_sc_hd__mux2_1 _11279_ (.A0(_05518_),
    .A1(\data_array.data1[10][49] ),
    .S(_05548_),
    .X(_03022_));
 sky130_fd_sc_hd__mux2_1 _11280_ (.A0(_05520_),
    .A1(\data_array.data1[10][50] ),
    .S(_05548_),
    .X(_03023_));
 sky130_fd_sc_hd__mux2_1 _11281_ (.A0(_05522_),
    .A1(\data_array.data1[10][51] ),
    .S(_05548_),
    .X(_03024_));
 sky130_fd_sc_hd__mux2_1 _11282_ (.A0(_05524_),
    .A1(\data_array.data1[10][52] ),
    .S(_05548_),
    .X(_03025_));
 sky130_fd_sc_hd__mux2_1 _11283_ (.A0(_05526_),
    .A1(\data_array.data1[10][53] ),
    .S(_05548_),
    .X(_03026_));
 sky130_fd_sc_hd__mux2_1 _11284_ (.A0(_05528_),
    .A1(\data_array.data1[10][54] ),
    .S(_05548_),
    .X(_03027_));
 sky130_fd_sc_hd__mux2_1 _11285_ (.A0(_05530_),
    .A1(\data_array.data1[10][55] ),
    .S(_05548_),
    .X(_03028_));
 sky130_fd_sc_hd__mux2_1 _11286_ (.A0(_05532_),
    .A1(\data_array.data1[10][56] ),
    .S(_05548_),
    .X(_03029_));
 sky130_fd_sc_hd__mux2_1 _11287_ (.A0(_05534_),
    .A1(\data_array.data1[10][57] ),
    .S(_05548_),
    .X(_03030_));
 sky130_fd_sc_hd__mux2_1 _11288_ (.A0(_05536_),
    .A1(\data_array.data1[10][58] ),
    .S(_05548_),
    .X(_03031_));
 sky130_fd_sc_hd__mux2_1 _11289_ (.A0(_05538_),
    .A1(\data_array.data1[10][59] ),
    .S(_05548_),
    .X(_03032_));
 sky130_fd_sc_hd__mux2_1 _11290_ (.A0(_05540_),
    .A1(\data_array.data1[10][60] ),
    .S(_05548_),
    .X(_03033_));
 sky130_fd_sc_hd__mux2_1 _11291_ (.A0(_05542_),
    .A1(\data_array.data1[10][61] ),
    .S(_05548_),
    .X(_03034_));
 sky130_fd_sc_hd__mux2_1 _11292_ (.A0(_05544_),
    .A1(\data_array.data1[10][62] ),
    .S(_05548_),
    .X(_03035_));
 sky130_fd_sc_hd__mux2_1 _11293_ (.A0(_05546_),
    .A1(\data_array.data1[10][63] ),
    .S(_05548_),
    .X(_03036_));
 sky130_fd_sc_hd__mux2_1 _11294_ (.A0(_05356_),
    .A1(\lru_array.lru_mem[13] ),
    .S(_05559_),
    .X(_03037_));
 sky130_fd_sc_hd__mux2_1 _11295_ (.A0(_05356_),
    .A1(\lru_array.lru_mem[14] ),
    .S(_05553_),
    .X(_03038_));
 sky130_fd_sc_hd__mux2_1 _11296_ (.A0(_05420_),
    .A1(\data_array.data1[7][0] ),
    .S(_05362_),
    .X(_03039_));
 sky130_fd_sc_hd__mux2_1 _11297_ (.A0(_05422_),
    .A1(\data_array.data1[7][1] ),
    .S(_05362_),
    .X(_03040_));
 sky130_fd_sc_hd__mux2_1 _11298_ (.A0(_05424_),
    .A1(\data_array.data1[7][2] ),
    .S(_05362_),
    .X(_03041_));
 sky130_fd_sc_hd__mux2_1 _11299_ (.A0(_05426_),
    .A1(\data_array.data1[7][3] ),
    .S(_05362_),
    .X(_03042_));
 sky130_fd_sc_hd__mux2_1 _11300_ (.A0(_05428_),
    .A1(\data_array.data1[7][4] ),
    .S(_05362_),
    .X(_03043_));
 sky130_fd_sc_hd__mux2_1 _11301_ (.A0(_05430_),
    .A1(\data_array.data1[7][5] ),
    .S(_05362_),
    .X(_03044_));
 sky130_fd_sc_hd__mux2_1 _11302_ (.A0(_05432_),
    .A1(\data_array.data1[7][6] ),
    .S(_05362_),
    .X(_03045_));
 sky130_fd_sc_hd__mux2_1 _11303_ (.A0(_05434_),
    .A1(\data_array.data1[7][7] ),
    .S(_05362_),
    .X(_03046_));
 sky130_fd_sc_hd__mux2_1 _11304_ (.A0(_05436_),
    .A1(\data_array.data1[7][8] ),
    .S(_05362_),
    .X(_03047_));
 sky130_fd_sc_hd__mux2_1 _11305_ (.A0(_05438_),
    .A1(\data_array.data1[7][9] ),
    .S(_05362_),
    .X(_03048_));
 sky130_fd_sc_hd__mux2_1 _11306_ (.A0(_05440_),
    .A1(\data_array.data1[7][10] ),
    .S(_05362_),
    .X(_03049_));
 sky130_fd_sc_hd__mux2_1 _11307_ (.A0(_05442_),
    .A1(\data_array.data1[7][11] ),
    .S(_05362_),
    .X(_03050_));
 sky130_fd_sc_hd__mux2_1 _11308_ (.A0(_05444_),
    .A1(\data_array.data1[7][12] ),
    .S(_05362_),
    .X(_03051_));
 sky130_fd_sc_hd__mux2_1 _11309_ (.A0(_05446_),
    .A1(\data_array.data1[7][13] ),
    .S(_05362_),
    .X(_03052_));
 sky130_fd_sc_hd__mux2_1 _11310_ (.A0(_05448_),
    .A1(\data_array.data1[7][14] ),
    .S(_05362_),
    .X(_03053_));
 sky130_fd_sc_hd__mux2_1 _11311_ (.A0(_05450_),
    .A1(\data_array.data1[7][15] ),
    .S(_05362_),
    .X(_03054_));
 sky130_fd_sc_hd__mux2_1 _11312_ (.A0(_05452_),
    .A1(\data_array.data1[7][16] ),
    .S(_05362_),
    .X(_03055_));
 sky130_fd_sc_hd__mux2_1 _11313_ (.A0(_05454_),
    .A1(\data_array.data1[7][17] ),
    .S(_05362_),
    .X(_03056_));
 sky130_fd_sc_hd__mux2_1 _11314_ (.A0(_05456_),
    .A1(\data_array.data1[7][18] ),
    .S(_05362_),
    .X(_03057_));
 sky130_fd_sc_hd__mux2_1 _11315_ (.A0(_05458_),
    .A1(\data_array.data1[7][19] ),
    .S(_05362_),
    .X(_03058_));
 sky130_fd_sc_hd__mux2_1 _11316_ (.A0(_05460_),
    .A1(\data_array.data1[7][20] ),
    .S(_05362_),
    .X(_03059_));
 sky130_fd_sc_hd__mux2_1 _11317_ (.A0(_05462_),
    .A1(\data_array.data1[7][21] ),
    .S(_05362_),
    .X(_03060_));
 sky130_fd_sc_hd__mux2_1 _11318_ (.A0(_05464_),
    .A1(\data_array.data1[7][22] ),
    .S(_05362_),
    .X(_03061_));
 sky130_fd_sc_hd__mux2_1 _11319_ (.A0(_05466_),
    .A1(\data_array.data1[7][23] ),
    .S(_05362_),
    .X(_03062_));
 sky130_fd_sc_hd__mux2_1 _11320_ (.A0(_05468_),
    .A1(\data_array.data1[7][24] ),
    .S(_05362_),
    .X(_03063_));
 sky130_fd_sc_hd__mux2_1 _11321_ (.A0(_05470_),
    .A1(\data_array.data1[7][25] ),
    .S(_05362_),
    .X(_03064_));
 sky130_fd_sc_hd__mux2_1 _11322_ (.A0(_05472_),
    .A1(\data_array.data1[7][26] ),
    .S(_05362_),
    .X(_03065_));
 sky130_fd_sc_hd__mux2_1 _11323_ (.A0(_05474_),
    .A1(\data_array.data1[7][27] ),
    .S(_05362_),
    .X(_03066_));
 sky130_fd_sc_hd__mux2_1 _11324_ (.A0(_05476_),
    .A1(\data_array.data1[7][28] ),
    .S(_05362_),
    .X(_03067_));
 sky130_fd_sc_hd__mux2_1 _11325_ (.A0(_05478_),
    .A1(\data_array.data1[7][29] ),
    .S(_05362_),
    .X(_03068_));
 sky130_fd_sc_hd__mux2_1 _11326_ (.A0(_05480_),
    .A1(\data_array.data1[7][30] ),
    .S(_05362_),
    .X(_03069_));
 sky130_fd_sc_hd__mux2_1 _11327_ (.A0(_05482_),
    .A1(\data_array.data1[7][31] ),
    .S(_05362_),
    .X(_03070_));
 sky130_fd_sc_hd__mux2_1 _11328_ (.A0(_05484_),
    .A1(\data_array.data1[7][32] ),
    .S(_05362_),
    .X(_03071_));
 sky130_fd_sc_hd__mux2_1 _11329_ (.A0(_05486_),
    .A1(\data_array.data1[7][33] ),
    .S(_05362_),
    .X(_03072_));
 sky130_fd_sc_hd__mux2_1 _11330_ (.A0(_05488_),
    .A1(\data_array.data1[7][34] ),
    .S(_05362_),
    .X(_03073_));
 sky130_fd_sc_hd__mux2_1 _11331_ (.A0(_05490_),
    .A1(\data_array.data1[7][35] ),
    .S(_05362_),
    .X(_03074_));
 sky130_fd_sc_hd__mux2_1 _11332_ (.A0(_05492_),
    .A1(\data_array.data1[7][36] ),
    .S(_05362_),
    .X(_03075_));
 sky130_fd_sc_hd__mux2_1 _11333_ (.A0(_05494_),
    .A1(\data_array.data1[7][37] ),
    .S(_05362_),
    .X(_03076_));
 sky130_fd_sc_hd__mux2_1 _11334_ (.A0(_05496_),
    .A1(\data_array.data1[7][38] ),
    .S(_05362_),
    .X(_03077_));
 sky130_fd_sc_hd__mux2_1 _11335_ (.A0(_05498_),
    .A1(\data_array.data1[7][39] ),
    .S(_05362_),
    .X(_03078_));
 sky130_fd_sc_hd__mux2_1 _11336_ (.A0(_05500_),
    .A1(\data_array.data1[7][40] ),
    .S(_05362_),
    .X(_03079_));
 sky130_fd_sc_hd__mux2_1 _11337_ (.A0(_05502_),
    .A1(\data_array.data1[7][41] ),
    .S(_05362_),
    .X(_03080_));
 sky130_fd_sc_hd__mux2_1 _11338_ (.A0(_05504_),
    .A1(\data_array.data1[7][42] ),
    .S(_05362_),
    .X(_03081_));
 sky130_fd_sc_hd__mux2_1 _11339_ (.A0(_05506_),
    .A1(\data_array.data1[7][43] ),
    .S(_05362_),
    .X(_03082_));
 sky130_fd_sc_hd__mux2_1 _11340_ (.A0(_05508_),
    .A1(\data_array.data1[7][44] ),
    .S(_05362_),
    .X(_03083_));
 sky130_fd_sc_hd__mux2_1 _11341_ (.A0(_05510_),
    .A1(\data_array.data1[7][45] ),
    .S(_05362_),
    .X(_03084_));
 sky130_fd_sc_hd__mux2_1 _11342_ (.A0(_05512_),
    .A1(\data_array.data1[7][46] ),
    .S(_05362_),
    .X(_03085_));
 sky130_fd_sc_hd__mux2_1 _11343_ (.A0(_05514_),
    .A1(\data_array.data1[7][47] ),
    .S(_05362_),
    .X(_03086_));
 sky130_fd_sc_hd__mux2_1 _11344_ (.A0(_05516_),
    .A1(\data_array.data1[7][48] ),
    .S(_05362_),
    .X(_03087_));
 sky130_fd_sc_hd__mux2_1 _11345_ (.A0(_05518_),
    .A1(\data_array.data1[7][49] ),
    .S(_05362_),
    .X(_03088_));
 sky130_fd_sc_hd__mux2_1 _11346_ (.A0(_05520_),
    .A1(\data_array.data1[7][50] ),
    .S(_05362_),
    .X(_03089_));
 sky130_fd_sc_hd__mux2_1 _11347_ (.A0(_05522_),
    .A1(\data_array.data1[7][51] ),
    .S(_05362_),
    .X(_03090_));
 sky130_fd_sc_hd__mux2_1 _11348_ (.A0(_05524_),
    .A1(\data_array.data1[7][52] ),
    .S(_05362_),
    .X(_03091_));
 sky130_fd_sc_hd__mux2_1 _11349_ (.A0(_05526_),
    .A1(\data_array.data1[7][53] ),
    .S(_05362_),
    .X(_03092_));
 sky130_fd_sc_hd__mux2_1 _11350_ (.A0(_05528_),
    .A1(\data_array.data1[7][54] ),
    .S(_05362_),
    .X(_03093_));
 sky130_fd_sc_hd__mux2_1 _11351_ (.A0(_05530_),
    .A1(\data_array.data1[7][55] ),
    .S(_05362_),
    .X(_03094_));
 sky130_fd_sc_hd__mux2_1 _11352_ (.A0(_05532_),
    .A1(\data_array.data1[7][56] ),
    .S(_05362_),
    .X(_03095_));
 sky130_fd_sc_hd__mux2_1 _11353_ (.A0(_05534_),
    .A1(\data_array.data1[7][57] ),
    .S(_05362_),
    .X(_03096_));
 sky130_fd_sc_hd__mux2_1 _11354_ (.A0(_05536_),
    .A1(\data_array.data1[7][58] ),
    .S(_05362_),
    .X(_03097_));
 sky130_fd_sc_hd__mux2_1 _11355_ (.A0(_05538_),
    .A1(\data_array.data1[7][59] ),
    .S(_05362_),
    .X(_03098_));
 sky130_fd_sc_hd__mux2_1 _11356_ (.A0(_05540_),
    .A1(\data_array.data1[7][60] ),
    .S(_05362_),
    .X(_03099_));
 sky130_fd_sc_hd__mux2_1 _11357_ (.A0(_05542_),
    .A1(\data_array.data1[7][61] ),
    .S(_05362_),
    .X(_03100_));
 sky130_fd_sc_hd__mux2_1 _11358_ (.A0(_05544_),
    .A1(\data_array.data1[7][62] ),
    .S(_05362_),
    .X(_03101_));
 sky130_fd_sc_hd__mux2_1 _11359_ (.A0(_05546_),
    .A1(\data_array.data1[7][63] ),
    .S(_05362_),
    .X(_03102_));
 sky130_fd_sc_hd__mux2_1 _11360_ (.A0(_05356_),
    .A1(\lru_array.lru_mem[9] ),
    .S(_05605_),
    .X(_03103_));
 sky130_fd_sc_hd__mux2_1 _11361_ (.A0(cpu_write),
    .A1(\tag_array.dirty0[15] ),
    .S(_05597_),
    .X(_03104_));
 sky130_fd_sc_hd__mux2_1 _11362_ (.A0(cpu_write),
    .A1(\tag_array.dirty0[1] ),
    .S(_05589_),
    .X(_03105_));
 sky130_fd_sc_hd__mux2_1 _11363_ (.A0(cpu_write),
    .A1(\tag_array.dirty0[2] ),
    .S(_05586_),
    .X(_03106_));
 sky130_fd_sc_hd__mux2_1 _11364_ (.A0(cpu_write),
    .A1(\tag_array.dirty0[3] ),
    .S(_05585_),
    .X(_03107_));
 sky130_fd_sc_hd__mux2_1 _11365_ (.A0(cpu_write),
    .A1(\tag_array.dirty0[4] ),
    .S(_05582_),
    .X(_03108_));
 sky130_fd_sc_hd__mux2_1 _11366_ (.A0(cpu_write),
    .A1(\tag_array.dirty0[5] ),
    .S(_05579_),
    .X(_03109_));
 sky130_fd_sc_hd__mux2_1 _11367_ (.A0(cpu_write),
    .A1(\tag_array.dirty0[6] ),
    .S(_05576_),
    .X(_03110_));
 sky130_fd_sc_hd__mux2_1 _11368_ (.A0(cpu_write),
    .A1(\tag_array.dirty0[7] ),
    .S(_05573_),
    .X(_03111_));
 sky130_fd_sc_hd__mux2_1 _11369_ (.A0(cpu_write),
    .A1(\tag_array.dirty0[8] ),
    .S(_05571_),
    .X(_03112_));
 sky130_fd_sc_hd__mux2_1 _11370_ (.A0(cpu_write),
    .A1(\tag_array.dirty0[0] ),
    .S(_05569_),
    .X(_03113_));
 sky130_fd_sc_hd__mux2_1 _11371_ (.A0(cpu_write),
    .A1(\tag_array.dirty0[10] ),
    .S(_05567_),
    .X(_03114_));
 sky130_fd_sc_hd__mux2_1 _11372_ (.A0(cpu_write),
    .A1(\tag_array.dirty0[11] ),
    .S(_05565_),
    .X(_03115_));
 sky130_fd_sc_hd__mux2_1 _11373_ (.A0(cpu_write),
    .A1(\tag_array.dirty0[12] ),
    .S(_05563_),
    .X(_03116_));
 sky130_fd_sc_hd__mux2_1 _11374_ (.A0(cpu_write),
    .A1(\tag_array.dirty0[13] ),
    .S(_05560_),
    .X(_03117_));
 sky130_fd_sc_hd__mux2_1 _11375_ (.A0(_05356_),
    .A1(\lru_array.lru_mem[3] ),
    .S(_05584_),
    .X(_03118_));
 sky130_fd_sc_hd__mux2_1 _11376_ (.A0(cpu_write),
    .A1(\tag_array.dirty0[14] ),
    .S(_05555_),
    .X(_03119_));
 sky130_fd_sc_hd__mux2_1 _11377_ (.A0(_05356_),
    .A1(\lru_array.lru_mem[12] ),
    .S(_05562_),
    .X(_03120_));
 sky130_fd_sc_hd__mux2_1 _11378_ (.A0(_05356_),
    .A1(\lru_array.lru_mem[4] ),
    .S(_05581_),
    .X(_03121_));
 sky130_fd_sc_hd__mux2_1 _11379_ (.A0(_05356_),
    .A1(\lru_array.lru_mem[5] ),
    .S(_05578_),
    .X(_03122_));
 sky130_fd_sc_hd__inv_2 _11380_ (.A(reset),
    .Y(_00190_));
 sky130_fd_sc_hd__inv_2 _11381_ (.A(reset),
    .Y(_00191_));
 sky130_fd_sc_hd__inv_2 _11382_ (.A(reset),
    .Y(_00192_));
 sky130_fd_sc_hd__inv_2 _11383_ (.A(reset),
    .Y(_00193_));
 sky130_fd_sc_hd__inv_2 _11384_ (.A(reset),
    .Y(_00194_));
 sky130_fd_sc_hd__dfxtp_2 _11385_ (.CLK(clk),
    .D(_00195_),
    .Q(\lru_array.lru_mem[2] ));
 sky130_fd_sc_hd__dfxtp_2 _11386_ (.CLK(clk),
    .D(_00196_),
    .Q(\tag_array.tag1[7][0] ));
 sky130_fd_sc_hd__dfxtp_2 _11387_ (.CLK(clk),
    .D(_00197_),
    .Q(\tag_array.tag1[7][1] ));
 sky130_fd_sc_hd__dfxtp_2 _11388_ (.CLK(clk),
    .D(_00198_),
    .Q(\tag_array.tag1[7][2] ));
 sky130_fd_sc_hd__dfxtp_2 _11389_ (.CLK(clk),
    .D(_00199_),
    .Q(\tag_array.tag1[7][3] ));
 sky130_fd_sc_hd__dfxtp_2 _11390_ (.CLK(clk),
    .D(_00200_),
    .Q(\tag_array.tag1[7][4] ));
 sky130_fd_sc_hd__dfxtp_2 _11391_ (.CLK(clk),
    .D(_00201_),
    .Q(\tag_array.tag1[7][5] ));
 sky130_fd_sc_hd__dfxtp_2 _11392_ (.CLK(clk),
    .D(_00202_),
    .Q(\tag_array.tag1[7][6] ));
 sky130_fd_sc_hd__dfxtp_2 _11393_ (.CLK(clk),
    .D(_00203_),
    .Q(\tag_array.tag1[7][7] ));
 sky130_fd_sc_hd__dfxtp_2 _11394_ (.CLK(clk),
    .D(_00204_),
    .Q(\tag_array.tag1[7][8] ));
 sky130_fd_sc_hd__dfxtp_2 _11395_ (.CLK(clk),
    .D(_00205_),
    .Q(\tag_array.tag1[7][9] ));
 sky130_fd_sc_hd__dfxtp_2 _11396_ (.CLK(clk),
    .D(_00206_),
    .Q(\tag_array.tag1[7][10] ));
 sky130_fd_sc_hd__dfxtp_2 _11397_ (.CLK(clk),
    .D(_00207_),
    .Q(\tag_array.tag1[7][11] ));
 sky130_fd_sc_hd__dfxtp_2 _11398_ (.CLK(clk),
    .D(_00208_),
    .Q(\tag_array.tag1[7][12] ));
 sky130_fd_sc_hd__dfxtp_2 _11399_ (.CLK(clk),
    .D(_00209_),
    .Q(\tag_array.tag1[7][13] ));
 sky130_fd_sc_hd__dfxtp_2 _11400_ (.CLK(clk),
    .D(_00210_),
    .Q(\tag_array.tag1[7][14] ));
 sky130_fd_sc_hd__dfxtp_2 _11401_ (.CLK(clk),
    .D(_00211_),
    .Q(\tag_array.tag1[7][15] ));
 sky130_fd_sc_hd__dfxtp_2 _11402_ (.CLK(clk),
    .D(_00212_),
    .Q(\tag_array.tag1[7][16] ));
 sky130_fd_sc_hd__dfxtp_2 _11403_ (.CLK(clk),
    .D(_00213_),
    .Q(\tag_array.tag1[7][17] ));
 sky130_fd_sc_hd__dfxtp_2 _11404_ (.CLK(clk),
    .D(_00214_),
    .Q(\tag_array.tag1[7][18] ));
 sky130_fd_sc_hd__dfxtp_2 _11405_ (.CLK(clk),
    .D(_00215_),
    .Q(\tag_array.tag1[7][19] ));
 sky130_fd_sc_hd__dfxtp_2 _11406_ (.CLK(clk),
    .D(_00216_),
    .Q(\tag_array.tag1[7][20] ));
 sky130_fd_sc_hd__dfxtp_2 _11407_ (.CLK(clk),
    .D(_00217_),
    .Q(\tag_array.tag1[7][21] ));
 sky130_fd_sc_hd__dfxtp_2 _11408_ (.CLK(clk),
    .D(_00218_),
    .Q(\tag_array.tag1[7][22] ));
 sky130_fd_sc_hd__dfxtp_2 _11409_ (.CLK(clk),
    .D(_00219_),
    .Q(\tag_array.tag1[7][23] ));
 sky130_fd_sc_hd__dfxtp_2 _11410_ (.CLK(clk),
    .D(_00220_),
    .Q(\tag_array.tag1[7][24] ));
 sky130_fd_sc_hd__dfxtp_2 _11411_ (.CLK(clk),
    .D(_00221_),
    .Q(\data_array.data0[0][0] ));
 sky130_fd_sc_hd__dfxtp_2 _11412_ (.CLK(clk),
    .D(_00222_),
    .Q(\data_array.data0[0][1] ));
 sky130_fd_sc_hd__dfxtp_2 _11413_ (.CLK(clk),
    .D(_00223_),
    .Q(\data_array.data0[0][2] ));
 sky130_fd_sc_hd__dfxtp_2 _11414_ (.CLK(clk),
    .D(_00224_),
    .Q(\data_array.data0[0][3] ));
 sky130_fd_sc_hd__dfxtp_2 _11415_ (.CLK(clk),
    .D(_00225_),
    .Q(\data_array.data0[0][4] ));
 sky130_fd_sc_hd__dfxtp_2 _11416_ (.CLK(clk),
    .D(_00226_),
    .Q(\data_array.data0[0][5] ));
 sky130_fd_sc_hd__dfxtp_2 _11417_ (.CLK(clk),
    .D(_00227_),
    .Q(\data_array.data0[0][6] ));
 sky130_fd_sc_hd__dfxtp_2 _11418_ (.CLK(clk),
    .D(_00228_),
    .Q(\data_array.data0[0][7] ));
 sky130_fd_sc_hd__dfxtp_2 _11419_ (.CLK(clk),
    .D(_00229_),
    .Q(\data_array.data0[0][8] ));
 sky130_fd_sc_hd__dfxtp_2 _11420_ (.CLK(clk),
    .D(_00230_),
    .Q(\data_array.data0[0][9] ));
 sky130_fd_sc_hd__dfxtp_2 _11421_ (.CLK(clk),
    .D(_00231_),
    .Q(\data_array.data0[0][10] ));
 sky130_fd_sc_hd__dfxtp_2 _11422_ (.CLK(clk),
    .D(_00232_),
    .Q(\data_array.data0[0][11] ));
 sky130_fd_sc_hd__dfxtp_2 _11423_ (.CLK(clk),
    .D(_00233_),
    .Q(\data_array.data0[0][12] ));
 sky130_fd_sc_hd__dfxtp_2 _11424_ (.CLK(clk),
    .D(_00234_),
    .Q(\data_array.data0[0][13] ));
 sky130_fd_sc_hd__dfxtp_2 _11425_ (.CLK(clk),
    .D(_00235_),
    .Q(\data_array.data0[0][14] ));
 sky130_fd_sc_hd__dfxtp_2 _11426_ (.CLK(clk),
    .D(_00236_),
    .Q(\data_array.data0[0][15] ));
 sky130_fd_sc_hd__dfxtp_2 _11427_ (.CLK(clk),
    .D(_00237_),
    .Q(\data_array.data0[0][16] ));
 sky130_fd_sc_hd__dfxtp_2 _11428_ (.CLK(clk),
    .D(_00238_),
    .Q(\data_array.data0[0][17] ));
 sky130_fd_sc_hd__dfxtp_2 _11429_ (.CLK(clk),
    .D(_00239_),
    .Q(\data_array.data0[0][18] ));
 sky130_fd_sc_hd__dfxtp_2 _11430_ (.CLK(clk),
    .D(_00240_),
    .Q(\data_array.data0[0][19] ));
 sky130_fd_sc_hd__dfxtp_2 _11431_ (.CLK(clk),
    .D(_00241_),
    .Q(\data_array.data0[0][20] ));
 sky130_fd_sc_hd__dfxtp_2 _11432_ (.CLK(clk),
    .D(_00242_),
    .Q(\data_array.data0[0][21] ));
 sky130_fd_sc_hd__dfxtp_2 _11433_ (.CLK(clk),
    .D(_00243_),
    .Q(\data_array.data0[0][22] ));
 sky130_fd_sc_hd__dfxtp_2 _11434_ (.CLK(clk),
    .D(_00244_),
    .Q(\data_array.data0[0][23] ));
 sky130_fd_sc_hd__dfxtp_2 _11435_ (.CLK(clk),
    .D(_00245_),
    .Q(\data_array.data0[0][24] ));
 sky130_fd_sc_hd__dfxtp_2 _11436_ (.CLK(clk),
    .D(_00246_),
    .Q(\data_array.data0[0][25] ));
 sky130_fd_sc_hd__dfxtp_2 _11437_ (.CLK(clk),
    .D(_00247_),
    .Q(\data_array.data0[0][26] ));
 sky130_fd_sc_hd__dfxtp_2 _11438_ (.CLK(clk),
    .D(_00248_),
    .Q(\data_array.data0[0][27] ));
 sky130_fd_sc_hd__dfxtp_2 _11439_ (.CLK(clk),
    .D(_00249_),
    .Q(\data_array.data0[0][28] ));
 sky130_fd_sc_hd__dfxtp_2 _11440_ (.CLK(clk),
    .D(_00250_),
    .Q(\data_array.data0[0][29] ));
 sky130_fd_sc_hd__dfxtp_2 _11441_ (.CLK(clk),
    .D(_00251_),
    .Q(\data_array.data0[0][30] ));
 sky130_fd_sc_hd__dfxtp_2 _11442_ (.CLK(clk),
    .D(_00252_),
    .Q(\data_array.data0[0][31] ));
 sky130_fd_sc_hd__dfxtp_2 _11443_ (.CLK(clk),
    .D(_00253_),
    .Q(\data_array.data0[0][32] ));
 sky130_fd_sc_hd__dfxtp_2 _11444_ (.CLK(clk),
    .D(_00254_),
    .Q(\data_array.data0[0][33] ));
 sky130_fd_sc_hd__dfxtp_2 _11445_ (.CLK(clk),
    .D(_00255_),
    .Q(\data_array.data0[0][34] ));
 sky130_fd_sc_hd__dfxtp_2 _11446_ (.CLK(clk),
    .D(_00256_),
    .Q(\data_array.data0[0][35] ));
 sky130_fd_sc_hd__dfxtp_2 _11447_ (.CLK(clk),
    .D(_00257_),
    .Q(\data_array.data0[0][36] ));
 sky130_fd_sc_hd__dfxtp_2 _11448_ (.CLK(clk),
    .D(_00258_),
    .Q(\data_array.data0[0][37] ));
 sky130_fd_sc_hd__dfxtp_2 _11449_ (.CLK(clk),
    .D(_00259_),
    .Q(\data_array.data0[0][38] ));
 sky130_fd_sc_hd__dfxtp_2 _11450_ (.CLK(clk),
    .D(_00260_),
    .Q(\data_array.data0[0][39] ));
 sky130_fd_sc_hd__dfxtp_2 _11451_ (.CLK(clk),
    .D(_00261_),
    .Q(\data_array.data0[0][40] ));
 sky130_fd_sc_hd__dfxtp_2 _11452_ (.CLK(clk),
    .D(_00262_),
    .Q(\data_array.data0[0][41] ));
 sky130_fd_sc_hd__dfxtp_2 _11453_ (.CLK(clk),
    .D(_00263_),
    .Q(\data_array.data0[0][42] ));
 sky130_fd_sc_hd__dfxtp_2 _11454_ (.CLK(clk),
    .D(_00264_),
    .Q(\data_array.data0[0][43] ));
 sky130_fd_sc_hd__dfxtp_2 _11455_ (.CLK(clk),
    .D(_00265_),
    .Q(\data_array.data0[0][44] ));
 sky130_fd_sc_hd__dfxtp_2 _11456_ (.CLK(clk),
    .D(_00266_),
    .Q(\data_array.data0[0][45] ));
 sky130_fd_sc_hd__dfxtp_2 _11457_ (.CLK(clk),
    .D(_00267_),
    .Q(\data_array.data0[0][46] ));
 sky130_fd_sc_hd__dfxtp_2 _11458_ (.CLK(clk),
    .D(_00268_),
    .Q(\data_array.data0[0][47] ));
 sky130_fd_sc_hd__dfxtp_2 _11459_ (.CLK(clk),
    .D(_00269_),
    .Q(\data_array.data0[0][48] ));
 sky130_fd_sc_hd__dfxtp_2 _11460_ (.CLK(clk),
    .D(_00270_),
    .Q(\data_array.data0[0][49] ));
 sky130_fd_sc_hd__dfxtp_2 _11461_ (.CLK(clk),
    .D(_00271_),
    .Q(\data_array.data0[0][50] ));
 sky130_fd_sc_hd__dfxtp_2 _11462_ (.CLK(clk),
    .D(_00272_),
    .Q(\data_array.data0[0][51] ));
 sky130_fd_sc_hd__dfxtp_2 _11463_ (.CLK(clk),
    .D(_00273_),
    .Q(\data_array.data0[0][52] ));
 sky130_fd_sc_hd__dfxtp_2 _11464_ (.CLK(clk),
    .D(_00274_),
    .Q(\data_array.data0[0][53] ));
 sky130_fd_sc_hd__dfxtp_2 _11465_ (.CLK(clk),
    .D(_00275_),
    .Q(\data_array.data0[0][54] ));
 sky130_fd_sc_hd__dfxtp_2 _11466_ (.CLK(clk),
    .D(_00276_),
    .Q(\data_array.data0[0][55] ));
 sky130_fd_sc_hd__dfxtp_2 _11467_ (.CLK(clk),
    .D(_00277_),
    .Q(\data_array.data0[0][56] ));
 sky130_fd_sc_hd__dfxtp_2 _11468_ (.CLK(clk),
    .D(_00278_),
    .Q(\data_array.data0[0][57] ));
 sky130_fd_sc_hd__dfxtp_2 _11469_ (.CLK(clk),
    .D(_00279_),
    .Q(\data_array.data0[0][58] ));
 sky130_fd_sc_hd__dfxtp_2 _11470_ (.CLK(clk),
    .D(_00280_),
    .Q(\data_array.data0[0][59] ));
 sky130_fd_sc_hd__dfxtp_2 _11471_ (.CLK(clk),
    .D(_00281_),
    .Q(\data_array.data0[0][60] ));
 sky130_fd_sc_hd__dfxtp_2 _11472_ (.CLK(clk),
    .D(_00282_),
    .Q(\data_array.data0[0][61] ));
 sky130_fd_sc_hd__dfxtp_2 _11473_ (.CLK(clk),
    .D(_00283_),
    .Q(\data_array.data0[0][62] ));
 sky130_fd_sc_hd__dfxtp_2 _11474_ (.CLK(clk),
    .D(_00284_),
    .Q(\data_array.data0[0][63] ));
 sky130_fd_sc_hd__dfxtp_2 _11475_ (.CLK(clk),
    .D(_00285_),
    .Q(\tag_array.valid1[10] ));
 sky130_fd_sc_hd__dfxtp_2 _11476_ (.CLK(clk),
    .D(_00286_),
    .Q(\tag_array.valid1[0] ));
 sky130_fd_sc_hd__dfxtp_2 _11477_ (.CLK(clk),
    .D(_00287_),
    .Q(\tag_array.valid1[11] ));
 sky130_fd_sc_hd__dfxtp_2 _11478_ (.CLK(clk),
    .D(_00181_),
    .Q(\fsm.valid0 ));
 sky130_fd_sc_hd__dfxtp_2 _11479_ (.CLK(clk),
    .D(_00288_),
    .Q(\tag_array.valid0[14] ));
 sky130_fd_sc_hd__dfxtp_2 _11480_ (.CLK(clk),
    .D(_00289_),
    .Q(\tag_array.valid1[8] ));
 sky130_fd_sc_hd__dfxtp_2 _11481_ (.CLK(clk),
    .D(_00290_),
    .Q(\tag_array.valid0[13] ));
 sky130_fd_sc_hd__dfxtp_2 _11482_ (.CLK(clk),
    .D(_00291_),
    .Q(\tag_array.valid1[7] ));
 sky130_fd_sc_hd__dfxtp_2 _11483_ (.CLK(clk),
    .D(_00292_),
    .Q(\tag_array.valid0[12] ));
 sky130_fd_sc_hd__dfxtp_2 _11484_ (.CLK(clk),
    .D(_00293_),
    .Q(\tag_array.valid0[11] ));
 sky130_fd_sc_hd__dfxtp_2 _11485_ (.CLK(clk),
    .D(_00294_),
    .Q(\tag_array.valid0[10] ));
 sky130_fd_sc_hd__dfxtp_2 _11486_ (.CLK(clk),
    .D(_00295_),
    .Q(\tag_array.valid0[0] ));
 sky130_fd_sc_hd__dfxtp_2 _11487_ (.CLK(clk),
    .D(_00296_),
    .Q(\tag_array.valid0[8] ));
 sky130_fd_sc_hd__dfxtp_2 _11488_ (.CLK(clk),
    .D(_00297_),
    .Q(\tag_array.valid0[7] ));
 sky130_fd_sc_hd__dfxtp_2 _11489_ (.CLK(clk),
    .D(_00298_),
    .Q(\tag_array.valid0[6] ));
 sky130_fd_sc_hd__dfxtp_2 _11490_ (.CLK(clk),
    .D(_00299_),
    .Q(\tag_array.valid0[5] ));
 sky130_fd_sc_hd__dfxtp_2 _11491_ (.CLK(clk),
    .D(_00300_),
    .Q(\tag_array.valid0[4] ));
 sky130_fd_sc_hd__dfxtp_2 _11492_ (.CLK(clk),
    .D(_00301_),
    .Q(\tag_array.valid0[3] ));
 sky130_fd_sc_hd__dfxtp_2 _11493_ (.CLK(clk),
    .D(_00302_),
    .Q(\tag_array.valid0[2] ));
 sky130_fd_sc_hd__dfxtp_2 _11494_ (.CLK(clk),
    .D(_00303_),
    .Q(\tag_array.valid0[1] ));
 sky130_fd_sc_hd__dfxtp_2 _11495_ (.CLK(clk),
    .D(_00304_),
    .Q(\tag_array.valid1[9] ));
 sky130_fd_sc_hd__dfxtp_2 _11496_ (.CLK(clk),
    .D(_00182_),
    .Q(\fsm.valid1 ));
 sky130_fd_sc_hd__dfxtp_2 _11497_ (.CLK(clk),
    .D(_00305_),
    .Q(\tag_array.valid1[14] ));
 sky130_fd_sc_hd__dfxtp_2 _11498_ (.CLK(clk),
    .D(_00306_),
    .Q(\tag_array.valid1[13] ));
 sky130_fd_sc_hd__dfxtp_2 _11499_ (.CLK(clk),
    .D(_00307_),
    .Q(\tag_array.valid1[12] ));
 sky130_fd_sc_hd__dfxtp_2 _11500_ (.CLK(clk),
    .D(_00308_),
    .Q(\tag_array.valid0[15] ));
 sky130_fd_sc_hd__dfxtp_2 _11501_ (.CLK(clk),
    .D(_00309_),
    .Q(\tag_array.tag1[9][0] ));
 sky130_fd_sc_hd__dfxtp_2 _11502_ (.CLK(clk),
    .D(_00310_),
    .Q(\tag_array.tag1[9][1] ));
 sky130_fd_sc_hd__dfxtp_2 _11503_ (.CLK(clk),
    .D(_00311_),
    .Q(\tag_array.tag1[9][2] ));
 sky130_fd_sc_hd__dfxtp_2 _11504_ (.CLK(clk),
    .D(_00312_),
    .Q(\tag_array.tag1[9][3] ));
 sky130_fd_sc_hd__dfxtp_2 _11505_ (.CLK(clk),
    .D(_00313_),
    .Q(\tag_array.tag1[9][4] ));
 sky130_fd_sc_hd__dfxtp_2 _11506_ (.CLK(clk),
    .D(_00314_),
    .Q(\tag_array.tag1[9][5] ));
 sky130_fd_sc_hd__dfxtp_2 _11507_ (.CLK(clk),
    .D(_00315_),
    .Q(\tag_array.tag1[9][6] ));
 sky130_fd_sc_hd__dfxtp_2 _11508_ (.CLK(clk),
    .D(_00316_),
    .Q(\tag_array.tag1[9][7] ));
 sky130_fd_sc_hd__dfxtp_2 _11509_ (.CLK(clk),
    .D(_00317_),
    .Q(\tag_array.tag1[9][8] ));
 sky130_fd_sc_hd__dfxtp_2 _11510_ (.CLK(clk),
    .D(_00318_),
    .Q(\tag_array.tag1[9][9] ));
 sky130_fd_sc_hd__dfxtp_2 _11511_ (.CLK(clk),
    .D(_00319_),
    .Q(\tag_array.tag1[9][10] ));
 sky130_fd_sc_hd__dfxtp_2 _11512_ (.CLK(clk),
    .D(_00320_),
    .Q(\tag_array.tag1[9][11] ));
 sky130_fd_sc_hd__dfxtp_2 _11513_ (.CLK(clk),
    .D(_00321_),
    .Q(\tag_array.tag1[9][12] ));
 sky130_fd_sc_hd__dfxtp_2 _11514_ (.CLK(clk),
    .D(_00322_),
    .Q(\tag_array.tag1[9][13] ));
 sky130_fd_sc_hd__dfxtp_2 _11515_ (.CLK(clk),
    .D(_00323_),
    .Q(\tag_array.tag1[9][14] ));
 sky130_fd_sc_hd__dfxtp_2 _11516_ (.CLK(clk),
    .D(_00324_),
    .Q(\tag_array.tag1[9][15] ));
 sky130_fd_sc_hd__dfxtp_2 _11517_ (.CLK(clk),
    .D(_00325_),
    .Q(\tag_array.tag1[9][16] ));
 sky130_fd_sc_hd__dfxtp_2 _11518_ (.CLK(clk),
    .D(_00326_),
    .Q(\tag_array.tag1[9][17] ));
 sky130_fd_sc_hd__dfxtp_2 _11519_ (.CLK(clk),
    .D(_00327_),
    .Q(\tag_array.tag1[9][18] ));
 sky130_fd_sc_hd__dfxtp_2 _11520_ (.CLK(clk),
    .D(_00328_),
    .Q(\tag_array.tag1[9][19] ));
 sky130_fd_sc_hd__dfxtp_2 _11521_ (.CLK(clk),
    .D(_00329_),
    .Q(\tag_array.tag1[9][20] ));
 sky130_fd_sc_hd__dfxtp_2 _11522_ (.CLK(clk),
    .D(_00330_),
    .Q(\tag_array.tag1[9][21] ));
 sky130_fd_sc_hd__dfxtp_2 _11523_ (.CLK(clk),
    .D(_00331_),
    .Q(\tag_array.tag1[9][22] ));
 sky130_fd_sc_hd__dfxtp_2 _11524_ (.CLK(clk),
    .D(_00332_),
    .Q(\tag_array.tag1[9][23] ));
 sky130_fd_sc_hd__dfxtp_2 _11525_ (.CLK(clk),
    .D(_00333_),
    .Q(\tag_array.tag1[9][24] ));
 sky130_fd_sc_hd__dfxtp_2 _11526_ (.CLK(clk),
    .D(_00334_),
    .Q(\tag_array.valid1[6] ));
 sky130_fd_sc_hd__dfxtp_2 _11527_ (.CLK(clk),
    .D(_00335_),
    .Q(\tag_array.valid1[5] ));
 sky130_fd_sc_hd__dfxtp_2 _11528_ (.CLK(clk),
    .D(_00336_),
    .Q(\tag_array.valid1[4] ));
 sky130_fd_sc_hd__dfxtp_2 _11529_ (.CLK(clk),
    .D(_00337_),
    .Q(\tag_array.valid1[3] ));
 sky130_fd_sc_hd__dfxtp_2 _11530_ (.CLK(clk),
    .D(_00338_),
    .Q(\tag_array.valid1[2] ));
 sky130_fd_sc_hd__dfxtp_2 _11531_ (.CLK(clk),
    .D(_00339_),
    .Q(\tag_array.valid1[1] ));
 sky130_fd_sc_hd__dfxtp_2 _11532_ (.CLK(clk),
    .D(_00340_),
    .Q(\tag_array.valid1[15] ));
 sky130_fd_sc_hd__dfxtp_2 _11533_ (.CLK(clk),
    .D(_00341_),
    .Q(\tag_array.valid0[9] ));
 sky130_fd_sc_hd__dfxtp_2 _11534_ (.CLK(clk),
    .D(_00342_),
    .Q(\tag_array.tag1[6][0] ));
 sky130_fd_sc_hd__dfxtp_2 _11535_ (.CLK(clk),
    .D(_00343_),
    .Q(\tag_array.tag1[6][1] ));
 sky130_fd_sc_hd__dfxtp_2 _11536_ (.CLK(clk),
    .D(_00344_),
    .Q(\tag_array.tag1[6][2] ));
 sky130_fd_sc_hd__dfxtp_2 _11537_ (.CLK(clk),
    .D(_00345_),
    .Q(\tag_array.tag1[6][3] ));
 sky130_fd_sc_hd__dfxtp_2 _11538_ (.CLK(clk),
    .D(_00346_),
    .Q(\tag_array.tag1[6][4] ));
 sky130_fd_sc_hd__dfxtp_2 _11539_ (.CLK(clk),
    .D(_00347_),
    .Q(\tag_array.tag1[6][5] ));
 sky130_fd_sc_hd__dfxtp_2 _11540_ (.CLK(clk),
    .D(_00348_),
    .Q(\tag_array.tag1[6][6] ));
 sky130_fd_sc_hd__dfxtp_2 _11541_ (.CLK(clk),
    .D(_00349_),
    .Q(\tag_array.tag1[6][7] ));
 sky130_fd_sc_hd__dfxtp_2 _11542_ (.CLK(clk),
    .D(_00350_),
    .Q(\tag_array.tag1[6][8] ));
 sky130_fd_sc_hd__dfxtp_2 _11543_ (.CLK(clk),
    .D(_00351_),
    .Q(\tag_array.tag1[6][9] ));
 sky130_fd_sc_hd__dfxtp_2 _11544_ (.CLK(clk),
    .D(_00352_),
    .Q(\tag_array.tag1[6][10] ));
 sky130_fd_sc_hd__dfxtp_2 _11545_ (.CLK(clk),
    .D(_00353_),
    .Q(\tag_array.tag1[6][11] ));
 sky130_fd_sc_hd__dfxtp_2 _11546_ (.CLK(clk),
    .D(_00354_),
    .Q(\tag_array.tag1[6][12] ));
 sky130_fd_sc_hd__dfxtp_2 _11547_ (.CLK(clk),
    .D(_00355_),
    .Q(\tag_array.tag1[6][13] ));
 sky130_fd_sc_hd__dfxtp_2 _11548_ (.CLK(clk),
    .D(_00356_),
    .Q(\tag_array.tag1[6][14] ));
 sky130_fd_sc_hd__dfxtp_2 _11549_ (.CLK(clk),
    .D(_00357_),
    .Q(\tag_array.tag1[6][15] ));
 sky130_fd_sc_hd__dfxtp_2 _11550_ (.CLK(clk),
    .D(_00358_),
    .Q(\tag_array.tag1[6][16] ));
 sky130_fd_sc_hd__dfxtp_2 _11551_ (.CLK(clk),
    .D(_00359_),
    .Q(\tag_array.tag1[6][17] ));
 sky130_fd_sc_hd__dfxtp_2 _11552_ (.CLK(clk),
    .D(_00360_),
    .Q(\tag_array.tag1[6][18] ));
 sky130_fd_sc_hd__dfxtp_2 _11553_ (.CLK(clk),
    .D(_00361_),
    .Q(\tag_array.tag1[6][19] ));
 sky130_fd_sc_hd__dfxtp_2 _11554_ (.CLK(clk),
    .D(_00362_),
    .Q(\tag_array.tag1[6][20] ));
 sky130_fd_sc_hd__dfxtp_2 _11555_ (.CLK(clk),
    .D(_00363_),
    .Q(\tag_array.tag1[6][21] ));
 sky130_fd_sc_hd__dfxtp_2 _11556_ (.CLK(clk),
    .D(_00364_),
    .Q(\tag_array.tag1[6][22] ));
 sky130_fd_sc_hd__dfxtp_2 _11557_ (.CLK(clk),
    .D(_00365_),
    .Q(\tag_array.tag1[6][23] ));
 sky130_fd_sc_hd__dfxtp_2 _11558_ (.CLK(clk),
    .D(_00366_),
    .Q(\tag_array.tag1[6][24] ));
 sky130_fd_sc_hd__dfxtp_2 _11559_ (.CLK(clk),
    .D(_00367_),
    .Q(\tag_array.tag1[5][0] ));
 sky130_fd_sc_hd__dfxtp_2 _11560_ (.CLK(clk),
    .D(_00368_),
    .Q(\tag_array.tag1[5][1] ));
 sky130_fd_sc_hd__dfxtp_2 _11561_ (.CLK(clk),
    .D(_00369_),
    .Q(\tag_array.tag1[5][2] ));
 sky130_fd_sc_hd__dfxtp_2 _11562_ (.CLK(clk),
    .D(_00370_),
    .Q(\tag_array.tag1[5][3] ));
 sky130_fd_sc_hd__dfxtp_2 _11563_ (.CLK(clk),
    .D(_00371_),
    .Q(\tag_array.tag1[5][4] ));
 sky130_fd_sc_hd__dfxtp_2 _11564_ (.CLK(clk),
    .D(_00372_),
    .Q(\tag_array.tag1[5][5] ));
 sky130_fd_sc_hd__dfxtp_2 _11565_ (.CLK(clk),
    .D(_00373_),
    .Q(\tag_array.tag1[5][6] ));
 sky130_fd_sc_hd__dfxtp_2 _11566_ (.CLK(clk),
    .D(_00374_),
    .Q(\tag_array.tag1[5][7] ));
 sky130_fd_sc_hd__dfxtp_2 _11567_ (.CLK(clk),
    .D(_00375_),
    .Q(\tag_array.tag1[5][8] ));
 sky130_fd_sc_hd__dfxtp_2 _11568_ (.CLK(clk),
    .D(_00376_),
    .Q(\tag_array.tag1[5][9] ));
 sky130_fd_sc_hd__dfxtp_2 _11569_ (.CLK(clk),
    .D(_00377_),
    .Q(\tag_array.tag1[5][10] ));
 sky130_fd_sc_hd__dfxtp_2 _11570_ (.CLK(clk),
    .D(_00378_),
    .Q(\tag_array.tag1[5][11] ));
 sky130_fd_sc_hd__dfxtp_2 _11571_ (.CLK(clk),
    .D(_00379_),
    .Q(\tag_array.tag1[5][12] ));
 sky130_fd_sc_hd__dfxtp_2 _11572_ (.CLK(clk),
    .D(_00380_),
    .Q(\tag_array.tag1[5][13] ));
 sky130_fd_sc_hd__dfxtp_2 _11573_ (.CLK(clk),
    .D(_00381_),
    .Q(\tag_array.tag1[5][14] ));
 sky130_fd_sc_hd__dfxtp_2 _11574_ (.CLK(clk),
    .D(_00382_),
    .Q(\tag_array.tag1[5][15] ));
 sky130_fd_sc_hd__dfxtp_2 _11575_ (.CLK(clk),
    .D(_00383_),
    .Q(\tag_array.tag1[5][16] ));
 sky130_fd_sc_hd__dfxtp_2 _11576_ (.CLK(clk),
    .D(_00384_),
    .Q(\tag_array.tag1[5][17] ));
 sky130_fd_sc_hd__dfxtp_2 _11577_ (.CLK(clk),
    .D(_00385_),
    .Q(\tag_array.tag1[5][18] ));
 sky130_fd_sc_hd__dfxtp_2 _11578_ (.CLK(clk),
    .D(_00386_),
    .Q(\tag_array.tag1[5][19] ));
 sky130_fd_sc_hd__dfxtp_2 _11579_ (.CLK(clk),
    .D(_00387_),
    .Q(\tag_array.tag1[5][20] ));
 sky130_fd_sc_hd__dfxtp_2 _11580_ (.CLK(clk),
    .D(_00388_),
    .Q(\tag_array.tag1[5][21] ));
 sky130_fd_sc_hd__dfxtp_2 _11581_ (.CLK(clk),
    .D(_00389_),
    .Q(\tag_array.tag1[5][22] ));
 sky130_fd_sc_hd__dfxtp_2 _11582_ (.CLK(clk),
    .D(_00390_),
    .Q(\tag_array.tag1[5][23] ));
 sky130_fd_sc_hd__dfxtp_2 _11583_ (.CLK(clk),
    .D(_00391_),
    .Q(\tag_array.tag1[5][24] ));
 sky130_fd_sc_hd__dfxtp_2 _11584_ (.CLK(clk),
    .D(_00392_),
    .Q(\tag_array.tag1[4][0] ));
 sky130_fd_sc_hd__dfxtp_2 _11585_ (.CLK(clk),
    .D(_00393_),
    .Q(\tag_array.tag1[4][1] ));
 sky130_fd_sc_hd__dfxtp_2 _11586_ (.CLK(clk),
    .D(_00394_),
    .Q(\tag_array.tag1[4][2] ));
 sky130_fd_sc_hd__dfxtp_2 _11587_ (.CLK(clk),
    .D(_00395_),
    .Q(\tag_array.tag1[4][3] ));
 sky130_fd_sc_hd__dfxtp_2 _11588_ (.CLK(clk),
    .D(_00396_),
    .Q(\tag_array.tag1[4][4] ));
 sky130_fd_sc_hd__dfxtp_2 _11589_ (.CLK(clk),
    .D(_00397_),
    .Q(\tag_array.tag1[4][5] ));
 sky130_fd_sc_hd__dfxtp_2 _11590_ (.CLK(clk),
    .D(_00398_),
    .Q(\tag_array.tag1[4][6] ));
 sky130_fd_sc_hd__dfxtp_2 _11591_ (.CLK(clk),
    .D(_00399_),
    .Q(\tag_array.tag1[4][7] ));
 sky130_fd_sc_hd__dfxtp_2 _11592_ (.CLK(clk),
    .D(_00400_),
    .Q(\tag_array.tag1[4][8] ));
 sky130_fd_sc_hd__dfxtp_2 _11593_ (.CLK(clk),
    .D(_00401_),
    .Q(\tag_array.tag1[4][9] ));
 sky130_fd_sc_hd__dfxtp_2 _11594_ (.CLK(clk),
    .D(_00402_),
    .Q(\tag_array.tag1[4][10] ));
 sky130_fd_sc_hd__dfxtp_2 _11595_ (.CLK(clk),
    .D(_00403_),
    .Q(\tag_array.tag1[4][11] ));
 sky130_fd_sc_hd__dfxtp_2 _11596_ (.CLK(clk),
    .D(_00404_),
    .Q(\tag_array.tag1[4][12] ));
 sky130_fd_sc_hd__dfxtp_2 _11597_ (.CLK(clk),
    .D(_00405_),
    .Q(\tag_array.tag1[4][13] ));
 sky130_fd_sc_hd__dfxtp_2 _11598_ (.CLK(clk),
    .D(_00406_),
    .Q(\tag_array.tag1[4][14] ));
 sky130_fd_sc_hd__dfxtp_2 _11599_ (.CLK(clk),
    .D(_00407_),
    .Q(\tag_array.tag1[4][15] ));
 sky130_fd_sc_hd__dfxtp_2 _11600_ (.CLK(clk),
    .D(_00408_),
    .Q(\tag_array.tag1[4][16] ));
 sky130_fd_sc_hd__dfxtp_2 _11601_ (.CLK(clk),
    .D(_00409_),
    .Q(\tag_array.tag1[4][17] ));
 sky130_fd_sc_hd__dfxtp_2 _11602_ (.CLK(clk),
    .D(_00410_),
    .Q(\tag_array.tag1[4][18] ));
 sky130_fd_sc_hd__dfxtp_2 _11603_ (.CLK(clk),
    .D(_00411_),
    .Q(\tag_array.tag1[4][19] ));
 sky130_fd_sc_hd__dfxtp_2 _11604_ (.CLK(clk),
    .D(_00412_),
    .Q(\tag_array.tag1[4][20] ));
 sky130_fd_sc_hd__dfxtp_2 _11605_ (.CLK(clk),
    .D(_00413_),
    .Q(\tag_array.tag1[4][21] ));
 sky130_fd_sc_hd__dfxtp_2 _11606_ (.CLK(clk),
    .D(_00414_),
    .Q(\tag_array.tag1[4][22] ));
 sky130_fd_sc_hd__dfxtp_2 _11607_ (.CLK(clk),
    .D(_00415_),
    .Q(\tag_array.tag1[4][23] ));
 sky130_fd_sc_hd__dfxtp_2 _11608_ (.CLK(clk),
    .D(_00416_),
    .Q(\tag_array.tag1[4][24] ));
 sky130_fd_sc_hd__dfxtp_2 _11609_ (.CLK(clk),
    .D(_00417_),
    .Q(\tag_array.tag1[3][0] ));
 sky130_fd_sc_hd__dfxtp_2 _11610_ (.CLK(clk),
    .D(_00418_),
    .Q(\tag_array.tag1[3][1] ));
 sky130_fd_sc_hd__dfxtp_2 _11611_ (.CLK(clk),
    .D(_00419_),
    .Q(\tag_array.tag1[3][2] ));
 sky130_fd_sc_hd__dfxtp_2 _11612_ (.CLK(clk),
    .D(_00420_),
    .Q(\tag_array.tag1[3][3] ));
 sky130_fd_sc_hd__dfxtp_2 _11613_ (.CLK(clk),
    .D(_00421_),
    .Q(\tag_array.tag1[3][4] ));
 sky130_fd_sc_hd__dfxtp_2 _11614_ (.CLK(clk),
    .D(_00422_),
    .Q(\tag_array.tag1[3][5] ));
 sky130_fd_sc_hd__dfxtp_2 _11615_ (.CLK(clk),
    .D(_00423_),
    .Q(\tag_array.tag1[3][6] ));
 sky130_fd_sc_hd__dfxtp_2 _11616_ (.CLK(clk),
    .D(_00424_),
    .Q(\tag_array.tag1[3][7] ));
 sky130_fd_sc_hd__dfxtp_2 _11617_ (.CLK(clk),
    .D(_00425_),
    .Q(\tag_array.tag1[3][8] ));
 sky130_fd_sc_hd__dfxtp_2 _11618_ (.CLK(clk),
    .D(_00426_),
    .Q(\tag_array.tag1[3][9] ));
 sky130_fd_sc_hd__dfxtp_2 _11619_ (.CLK(clk),
    .D(_00427_),
    .Q(\tag_array.tag1[3][10] ));
 sky130_fd_sc_hd__dfxtp_2 _11620_ (.CLK(clk),
    .D(_00428_),
    .Q(\tag_array.tag1[3][11] ));
 sky130_fd_sc_hd__dfxtp_2 _11621_ (.CLK(clk),
    .D(_00429_),
    .Q(\tag_array.tag1[3][12] ));
 sky130_fd_sc_hd__dfxtp_2 _11622_ (.CLK(clk),
    .D(_00430_),
    .Q(\tag_array.tag1[3][13] ));
 sky130_fd_sc_hd__dfxtp_2 _11623_ (.CLK(clk),
    .D(_00431_),
    .Q(\tag_array.tag1[3][14] ));
 sky130_fd_sc_hd__dfxtp_2 _11624_ (.CLK(clk),
    .D(_00432_),
    .Q(\tag_array.tag1[3][15] ));
 sky130_fd_sc_hd__dfxtp_2 _11625_ (.CLK(clk),
    .D(_00433_),
    .Q(\tag_array.tag1[3][16] ));
 sky130_fd_sc_hd__dfxtp_2 _11626_ (.CLK(clk),
    .D(_00434_),
    .Q(\tag_array.tag1[3][17] ));
 sky130_fd_sc_hd__dfxtp_2 _11627_ (.CLK(clk),
    .D(_00435_),
    .Q(\tag_array.tag1[3][18] ));
 sky130_fd_sc_hd__dfxtp_2 _11628_ (.CLK(clk),
    .D(_00436_),
    .Q(\tag_array.tag1[3][19] ));
 sky130_fd_sc_hd__dfxtp_2 _11629_ (.CLK(clk),
    .D(_00437_),
    .Q(\tag_array.tag1[3][20] ));
 sky130_fd_sc_hd__dfxtp_2 _11630_ (.CLK(clk),
    .D(_00438_),
    .Q(\tag_array.tag1[3][21] ));
 sky130_fd_sc_hd__dfxtp_2 _11631_ (.CLK(clk),
    .D(_00439_),
    .Q(\tag_array.tag1[3][22] ));
 sky130_fd_sc_hd__dfxtp_2 _11632_ (.CLK(clk),
    .D(_00440_),
    .Q(\tag_array.tag1[3][23] ));
 sky130_fd_sc_hd__dfxtp_2 _11633_ (.CLK(clk),
    .D(_00441_),
    .Q(\tag_array.tag1[3][24] ));
 sky130_fd_sc_hd__dfxtp_2 _11634_ (.CLK(clk),
    .D(_00442_),
    .Q(\tag_array.tag1[2][0] ));
 sky130_fd_sc_hd__dfxtp_2 _11635_ (.CLK(clk),
    .D(_00443_),
    .Q(\tag_array.tag1[2][1] ));
 sky130_fd_sc_hd__dfxtp_2 _11636_ (.CLK(clk),
    .D(_00444_),
    .Q(\tag_array.tag1[2][2] ));
 sky130_fd_sc_hd__dfxtp_2 _11637_ (.CLK(clk),
    .D(_00445_),
    .Q(\tag_array.tag1[2][3] ));
 sky130_fd_sc_hd__dfxtp_2 _11638_ (.CLK(clk),
    .D(_00446_),
    .Q(\tag_array.tag1[2][4] ));
 sky130_fd_sc_hd__dfxtp_2 _11639_ (.CLK(clk),
    .D(_00447_),
    .Q(\tag_array.tag1[2][5] ));
 sky130_fd_sc_hd__dfxtp_2 _11640_ (.CLK(clk),
    .D(_00448_),
    .Q(\tag_array.tag1[2][6] ));
 sky130_fd_sc_hd__dfxtp_2 _11641_ (.CLK(clk),
    .D(_00449_),
    .Q(\tag_array.tag1[2][7] ));
 sky130_fd_sc_hd__dfxtp_2 _11642_ (.CLK(clk),
    .D(_00450_),
    .Q(\tag_array.tag1[2][8] ));
 sky130_fd_sc_hd__dfxtp_2 _11643_ (.CLK(clk),
    .D(_00451_),
    .Q(\tag_array.tag1[2][9] ));
 sky130_fd_sc_hd__dfxtp_2 _11644_ (.CLK(clk),
    .D(_00452_),
    .Q(\tag_array.tag1[2][10] ));
 sky130_fd_sc_hd__dfxtp_2 _11645_ (.CLK(clk),
    .D(_00453_),
    .Q(\tag_array.tag1[2][11] ));
 sky130_fd_sc_hd__dfxtp_2 _11646_ (.CLK(clk),
    .D(_00454_),
    .Q(\tag_array.tag1[2][12] ));
 sky130_fd_sc_hd__dfxtp_2 _11647_ (.CLK(clk),
    .D(_00455_),
    .Q(\tag_array.tag1[2][13] ));
 sky130_fd_sc_hd__dfxtp_2 _11648_ (.CLK(clk),
    .D(_00456_),
    .Q(\tag_array.tag1[2][14] ));
 sky130_fd_sc_hd__dfxtp_2 _11649_ (.CLK(clk),
    .D(_00457_),
    .Q(\tag_array.tag1[2][15] ));
 sky130_fd_sc_hd__dfxtp_2 _11650_ (.CLK(clk),
    .D(_00458_),
    .Q(\tag_array.tag1[2][16] ));
 sky130_fd_sc_hd__dfxtp_2 _11651_ (.CLK(clk),
    .D(_00459_),
    .Q(\tag_array.tag1[2][17] ));
 sky130_fd_sc_hd__dfxtp_2 _11652_ (.CLK(clk),
    .D(_00460_),
    .Q(\tag_array.tag1[2][18] ));
 sky130_fd_sc_hd__dfxtp_2 _11653_ (.CLK(clk),
    .D(_00461_),
    .Q(\tag_array.tag1[2][19] ));
 sky130_fd_sc_hd__dfxtp_2 _11654_ (.CLK(clk),
    .D(_00462_),
    .Q(\tag_array.tag1[2][20] ));
 sky130_fd_sc_hd__dfxtp_2 _11655_ (.CLK(clk),
    .D(_00463_),
    .Q(\tag_array.tag1[2][21] ));
 sky130_fd_sc_hd__dfxtp_2 _11656_ (.CLK(clk),
    .D(_00464_),
    .Q(\tag_array.tag1[2][22] ));
 sky130_fd_sc_hd__dfxtp_2 _11657_ (.CLK(clk),
    .D(_00465_),
    .Q(\tag_array.tag1[2][23] ));
 sky130_fd_sc_hd__dfxtp_2 _11658_ (.CLK(clk),
    .D(_00466_),
    .Q(\tag_array.tag1[2][24] ));
 sky130_fd_sc_hd__dfxtp_2 _11659_ (.CLK(clk),
    .D(_00467_),
    .Q(\tag_array.tag1[1][0] ));
 sky130_fd_sc_hd__dfxtp_2 _11660_ (.CLK(clk),
    .D(_00468_),
    .Q(\tag_array.tag1[1][1] ));
 sky130_fd_sc_hd__dfxtp_2 _11661_ (.CLK(clk),
    .D(_00469_),
    .Q(\tag_array.tag1[1][2] ));
 sky130_fd_sc_hd__dfxtp_2 _11662_ (.CLK(clk),
    .D(_00470_),
    .Q(\tag_array.tag1[1][3] ));
 sky130_fd_sc_hd__dfxtp_2 _11663_ (.CLK(clk),
    .D(_00471_),
    .Q(\tag_array.tag1[1][4] ));
 sky130_fd_sc_hd__dfxtp_2 _11664_ (.CLK(clk),
    .D(_00472_),
    .Q(\tag_array.tag1[1][5] ));
 sky130_fd_sc_hd__dfxtp_2 _11665_ (.CLK(clk),
    .D(_00473_),
    .Q(\tag_array.tag1[1][6] ));
 sky130_fd_sc_hd__dfxtp_2 _11666_ (.CLK(clk),
    .D(_00474_),
    .Q(\tag_array.tag1[1][7] ));
 sky130_fd_sc_hd__dfxtp_2 _11667_ (.CLK(clk),
    .D(_00475_),
    .Q(\tag_array.tag1[1][8] ));
 sky130_fd_sc_hd__dfxtp_2 _11668_ (.CLK(clk),
    .D(_00476_),
    .Q(\tag_array.tag1[1][9] ));
 sky130_fd_sc_hd__dfxtp_2 _11669_ (.CLK(clk),
    .D(_00477_),
    .Q(\tag_array.tag1[1][10] ));
 sky130_fd_sc_hd__dfxtp_2 _11670_ (.CLK(clk),
    .D(_00478_),
    .Q(\tag_array.tag1[1][11] ));
 sky130_fd_sc_hd__dfxtp_2 _11671_ (.CLK(clk),
    .D(_00479_),
    .Q(\tag_array.tag1[1][12] ));
 sky130_fd_sc_hd__dfxtp_2 _11672_ (.CLK(clk),
    .D(_00480_),
    .Q(\tag_array.tag1[1][13] ));
 sky130_fd_sc_hd__dfxtp_2 _11673_ (.CLK(clk),
    .D(_00481_),
    .Q(\tag_array.tag1[1][14] ));
 sky130_fd_sc_hd__dfxtp_2 _11674_ (.CLK(clk),
    .D(_00482_),
    .Q(\tag_array.tag1[1][15] ));
 sky130_fd_sc_hd__dfxtp_2 _11675_ (.CLK(clk),
    .D(_00483_),
    .Q(\tag_array.tag1[1][16] ));
 sky130_fd_sc_hd__dfxtp_2 _11676_ (.CLK(clk),
    .D(_00484_),
    .Q(\tag_array.tag1[1][17] ));
 sky130_fd_sc_hd__dfxtp_2 _11677_ (.CLK(clk),
    .D(_00485_),
    .Q(\tag_array.tag1[1][18] ));
 sky130_fd_sc_hd__dfxtp_2 _11678_ (.CLK(clk),
    .D(_00486_),
    .Q(\tag_array.tag1[1][19] ));
 sky130_fd_sc_hd__dfxtp_2 _11679_ (.CLK(clk),
    .D(_00487_),
    .Q(\tag_array.tag1[1][20] ));
 sky130_fd_sc_hd__dfxtp_2 _11680_ (.CLK(clk),
    .D(_00488_),
    .Q(\tag_array.tag1[1][21] ));
 sky130_fd_sc_hd__dfxtp_2 _11681_ (.CLK(clk),
    .D(_00489_),
    .Q(\tag_array.tag1[1][22] ));
 sky130_fd_sc_hd__dfxtp_2 _11682_ (.CLK(clk),
    .D(_00490_),
    .Q(\tag_array.tag1[1][23] ));
 sky130_fd_sc_hd__dfxtp_2 _11683_ (.CLK(clk),
    .D(_00491_),
    .Q(\tag_array.tag1[1][24] ));
 sky130_fd_sc_hd__dfxtp_2 _11684_ (.CLK(clk),
    .D(_00492_),
    .Q(\tag_array.tag1[15][0] ));
 sky130_fd_sc_hd__dfxtp_2 _11685_ (.CLK(clk),
    .D(_00493_),
    .Q(\tag_array.tag1[15][1] ));
 sky130_fd_sc_hd__dfxtp_2 _11686_ (.CLK(clk),
    .D(_00494_),
    .Q(\tag_array.tag1[15][2] ));
 sky130_fd_sc_hd__dfxtp_2 _11687_ (.CLK(clk),
    .D(_00495_),
    .Q(\tag_array.tag1[15][3] ));
 sky130_fd_sc_hd__dfxtp_2 _11688_ (.CLK(clk),
    .D(_00496_),
    .Q(\tag_array.tag1[15][4] ));
 sky130_fd_sc_hd__dfxtp_2 _11689_ (.CLK(clk),
    .D(_00497_),
    .Q(\tag_array.tag1[15][5] ));
 sky130_fd_sc_hd__dfxtp_2 _11690_ (.CLK(clk),
    .D(_00498_),
    .Q(\tag_array.tag1[15][6] ));
 sky130_fd_sc_hd__dfxtp_2 _11691_ (.CLK(clk),
    .D(_00499_),
    .Q(\tag_array.tag1[15][7] ));
 sky130_fd_sc_hd__dfxtp_2 _11692_ (.CLK(clk),
    .D(_00500_),
    .Q(\tag_array.tag1[15][8] ));
 sky130_fd_sc_hd__dfxtp_2 _11693_ (.CLK(clk),
    .D(_00501_),
    .Q(\tag_array.tag1[15][9] ));
 sky130_fd_sc_hd__dfxtp_2 _11694_ (.CLK(clk),
    .D(_00502_),
    .Q(\tag_array.tag1[15][10] ));
 sky130_fd_sc_hd__dfxtp_2 _11695_ (.CLK(clk),
    .D(_00503_),
    .Q(\tag_array.tag1[15][11] ));
 sky130_fd_sc_hd__dfxtp_2 _11696_ (.CLK(clk),
    .D(_00504_),
    .Q(\tag_array.tag1[15][12] ));
 sky130_fd_sc_hd__dfxtp_2 _11697_ (.CLK(clk),
    .D(_00505_),
    .Q(\tag_array.tag1[15][13] ));
 sky130_fd_sc_hd__dfxtp_2 _11698_ (.CLK(clk),
    .D(_00506_),
    .Q(\tag_array.tag1[15][14] ));
 sky130_fd_sc_hd__dfxtp_2 _11699_ (.CLK(clk),
    .D(_00507_),
    .Q(\tag_array.tag1[15][15] ));
 sky130_fd_sc_hd__dfxtp_2 _11700_ (.CLK(clk),
    .D(_00508_),
    .Q(\tag_array.tag1[15][16] ));
 sky130_fd_sc_hd__dfxtp_2 _11701_ (.CLK(clk),
    .D(_00509_),
    .Q(\tag_array.tag1[15][17] ));
 sky130_fd_sc_hd__dfxtp_2 _11702_ (.CLK(clk),
    .D(_00510_),
    .Q(\tag_array.tag1[15][18] ));
 sky130_fd_sc_hd__dfxtp_2 _11703_ (.CLK(clk),
    .D(_00511_),
    .Q(\tag_array.tag1[15][19] ));
 sky130_fd_sc_hd__dfxtp_2 _11704_ (.CLK(clk),
    .D(_00512_),
    .Q(\tag_array.tag1[15][20] ));
 sky130_fd_sc_hd__dfxtp_2 _11705_ (.CLK(clk),
    .D(_00513_),
    .Q(\tag_array.tag1[15][21] ));
 sky130_fd_sc_hd__dfxtp_2 _11706_ (.CLK(clk),
    .D(_00514_),
    .Q(\tag_array.tag1[15][22] ));
 sky130_fd_sc_hd__dfxtp_2 _11707_ (.CLK(clk),
    .D(_00515_),
    .Q(\tag_array.tag1[15][23] ));
 sky130_fd_sc_hd__dfxtp_2 _11708_ (.CLK(clk),
    .D(_00516_),
    .Q(\tag_array.tag1[15][24] ));
 sky130_fd_sc_hd__dfxtp_2 _11709_ (.CLK(clk),
    .D(_00517_),
    .Q(\tag_array.tag0[9][0] ));
 sky130_fd_sc_hd__dfxtp_2 _11710_ (.CLK(clk),
    .D(_00518_),
    .Q(\tag_array.tag0[9][1] ));
 sky130_fd_sc_hd__dfxtp_2 _11711_ (.CLK(clk),
    .D(_00519_),
    .Q(\tag_array.tag0[9][2] ));
 sky130_fd_sc_hd__dfxtp_2 _11712_ (.CLK(clk),
    .D(_00520_),
    .Q(\tag_array.tag0[9][3] ));
 sky130_fd_sc_hd__dfxtp_2 _11713_ (.CLK(clk),
    .D(_00521_),
    .Q(\tag_array.tag0[9][4] ));
 sky130_fd_sc_hd__dfxtp_2 _11714_ (.CLK(clk),
    .D(_00522_),
    .Q(\tag_array.tag0[9][5] ));
 sky130_fd_sc_hd__dfxtp_2 _11715_ (.CLK(clk),
    .D(_00523_),
    .Q(\tag_array.tag0[9][6] ));
 sky130_fd_sc_hd__dfxtp_2 _11716_ (.CLK(clk),
    .D(_00524_),
    .Q(\tag_array.tag0[9][7] ));
 sky130_fd_sc_hd__dfxtp_2 _11717_ (.CLK(clk),
    .D(_00525_),
    .Q(\tag_array.tag0[9][8] ));
 sky130_fd_sc_hd__dfxtp_2 _11718_ (.CLK(clk),
    .D(_00526_),
    .Q(\tag_array.tag0[9][9] ));
 sky130_fd_sc_hd__dfxtp_2 _11719_ (.CLK(clk),
    .D(_00527_),
    .Q(\tag_array.tag0[9][10] ));
 sky130_fd_sc_hd__dfxtp_2 _11720_ (.CLK(clk),
    .D(_00528_),
    .Q(\tag_array.tag0[9][11] ));
 sky130_fd_sc_hd__dfxtp_2 _11721_ (.CLK(clk),
    .D(_00529_),
    .Q(\tag_array.tag0[9][12] ));
 sky130_fd_sc_hd__dfxtp_2 _11722_ (.CLK(clk),
    .D(_00530_),
    .Q(\tag_array.tag0[9][13] ));
 sky130_fd_sc_hd__dfxtp_2 _11723_ (.CLK(clk),
    .D(_00531_),
    .Q(\tag_array.tag0[9][14] ));
 sky130_fd_sc_hd__dfxtp_2 _11724_ (.CLK(clk),
    .D(_00532_),
    .Q(\tag_array.tag0[9][15] ));
 sky130_fd_sc_hd__dfxtp_2 _11725_ (.CLK(clk),
    .D(_00533_),
    .Q(\tag_array.tag0[9][16] ));
 sky130_fd_sc_hd__dfxtp_2 _11726_ (.CLK(clk),
    .D(_00534_),
    .Q(\tag_array.tag0[9][17] ));
 sky130_fd_sc_hd__dfxtp_2 _11727_ (.CLK(clk),
    .D(_00535_),
    .Q(\tag_array.tag0[9][18] ));
 sky130_fd_sc_hd__dfxtp_2 _11728_ (.CLK(clk),
    .D(_00536_),
    .Q(\tag_array.tag0[9][19] ));
 sky130_fd_sc_hd__dfxtp_2 _11729_ (.CLK(clk),
    .D(_00537_),
    .Q(\tag_array.tag0[9][20] ));
 sky130_fd_sc_hd__dfxtp_2 _11730_ (.CLK(clk),
    .D(_00538_),
    .Q(\tag_array.tag0[9][21] ));
 sky130_fd_sc_hd__dfxtp_2 _11731_ (.CLK(clk),
    .D(_00539_),
    .Q(\tag_array.tag0[9][22] ));
 sky130_fd_sc_hd__dfxtp_2 _11732_ (.CLK(clk),
    .D(_00540_),
    .Q(\tag_array.tag0[9][23] ));
 sky130_fd_sc_hd__dfxtp_2 _11733_ (.CLK(clk),
    .D(_00541_),
    .Q(\tag_array.tag0[9][24] ));
 sky130_fd_sc_hd__dfxtp_2 _11734_ (.CLK(clk),
    .D(_00542_),
    .Q(\data_array.data0[8][0] ));
 sky130_fd_sc_hd__dfxtp_2 _11735_ (.CLK(clk),
    .D(_00543_),
    .Q(\data_array.data0[8][1] ));
 sky130_fd_sc_hd__dfxtp_2 _11736_ (.CLK(clk),
    .D(_00544_),
    .Q(\data_array.data0[8][2] ));
 sky130_fd_sc_hd__dfxtp_2 _11737_ (.CLK(clk),
    .D(_00545_),
    .Q(\data_array.data0[8][3] ));
 sky130_fd_sc_hd__dfxtp_2 _11738_ (.CLK(clk),
    .D(_00546_),
    .Q(\data_array.data0[8][4] ));
 sky130_fd_sc_hd__dfxtp_2 _11739_ (.CLK(clk),
    .D(_00547_),
    .Q(\data_array.data0[8][5] ));
 sky130_fd_sc_hd__dfxtp_2 _11740_ (.CLK(clk),
    .D(_00548_),
    .Q(\data_array.data0[8][6] ));
 sky130_fd_sc_hd__dfxtp_2 _11741_ (.CLK(clk),
    .D(_00549_),
    .Q(\data_array.data0[8][7] ));
 sky130_fd_sc_hd__dfxtp_2 _11742_ (.CLK(clk),
    .D(_00550_),
    .Q(\data_array.data0[8][8] ));
 sky130_fd_sc_hd__dfxtp_2 _11743_ (.CLK(clk),
    .D(_00551_),
    .Q(\data_array.data0[8][9] ));
 sky130_fd_sc_hd__dfxtp_2 _11744_ (.CLK(clk),
    .D(_00552_),
    .Q(\data_array.data0[8][10] ));
 sky130_fd_sc_hd__dfxtp_2 _11745_ (.CLK(clk),
    .D(_00553_),
    .Q(\data_array.data0[8][11] ));
 sky130_fd_sc_hd__dfxtp_2 _11746_ (.CLK(clk),
    .D(_00554_),
    .Q(\data_array.data0[8][12] ));
 sky130_fd_sc_hd__dfxtp_2 _11747_ (.CLK(clk),
    .D(_00555_),
    .Q(\data_array.data0[8][13] ));
 sky130_fd_sc_hd__dfxtp_2 _11748_ (.CLK(clk),
    .D(_00556_),
    .Q(\data_array.data0[8][14] ));
 sky130_fd_sc_hd__dfxtp_2 _11749_ (.CLK(clk),
    .D(_00557_),
    .Q(\data_array.data0[8][15] ));
 sky130_fd_sc_hd__dfxtp_2 _11750_ (.CLK(clk),
    .D(_00558_),
    .Q(\data_array.data0[8][16] ));
 sky130_fd_sc_hd__dfxtp_2 _11751_ (.CLK(clk),
    .D(_00559_),
    .Q(\data_array.data0[8][17] ));
 sky130_fd_sc_hd__dfxtp_2 _11752_ (.CLK(clk),
    .D(_00560_),
    .Q(\data_array.data0[8][18] ));
 sky130_fd_sc_hd__dfxtp_2 _11753_ (.CLK(clk),
    .D(_00561_),
    .Q(\data_array.data0[8][19] ));
 sky130_fd_sc_hd__dfxtp_2 _11754_ (.CLK(clk),
    .D(_00562_),
    .Q(\data_array.data0[8][20] ));
 sky130_fd_sc_hd__dfxtp_2 _11755_ (.CLK(clk),
    .D(_00563_),
    .Q(\data_array.data0[8][21] ));
 sky130_fd_sc_hd__dfxtp_2 _11756_ (.CLK(clk),
    .D(_00564_),
    .Q(\data_array.data0[8][22] ));
 sky130_fd_sc_hd__dfxtp_2 _11757_ (.CLK(clk),
    .D(_00565_),
    .Q(\data_array.data0[8][23] ));
 sky130_fd_sc_hd__dfxtp_2 _11758_ (.CLK(clk),
    .D(_00566_),
    .Q(\data_array.data0[8][24] ));
 sky130_fd_sc_hd__dfxtp_2 _11759_ (.CLK(clk),
    .D(_00567_),
    .Q(\data_array.data0[8][25] ));
 sky130_fd_sc_hd__dfxtp_2 _11760_ (.CLK(clk),
    .D(_00568_),
    .Q(\data_array.data0[8][26] ));
 sky130_fd_sc_hd__dfxtp_2 _11761_ (.CLK(clk),
    .D(_00569_),
    .Q(\data_array.data0[8][27] ));
 sky130_fd_sc_hd__dfxtp_2 _11762_ (.CLK(clk),
    .D(_00570_),
    .Q(\data_array.data0[8][28] ));
 sky130_fd_sc_hd__dfxtp_2 _11763_ (.CLK(clk),
    .D(_00571_),
    .Q(\data_array.data0[8][29] ));
 sky130_fd_sc_hd__dfxtp_2 _11764_ (.CLK(clk),
    .D(_00572_),
    .Q(\data_array.data0[8][30] ));
 sky130_fd_sc_hd__dfxtp_2 _11765_ (.CLK(clk),
    .D(_00573_),
    .Q(\data_array.data0[8][31] ));
 sky130_fd_sc_hd__dfxtp_2 _11766_ (.CLK(clk),
    .D(_00574_),
    .Q(\data_array.data0[8][32] ));
 sky130_fd_sc_hd__dfxtp_2 _11767_ (.CLK(clk),
    .D(_00575_),
    .Q(\data_array.data0[8][33] ));
 sky130_fd_sc_hd__dfxtp_2 _11768_ (.CLK(clk),
    .D(_00576_),
    .Q(\data_array.data0[8][34] ));
 sky130_fd_sc_hd__dfxtp_2 _11769_ (.CLK(clk),
    .D(_00577_),
    .Q(\data_array.data0[8][35] ));
 sky130_fd_sc_hd__dfxtp_2 _11770_ (.CLK(clk),
    .D(_00578_),
    .Q(\data_array.data0[8][36] ));
 sky130_fd_sc_hd__dfxtp_2 _11771_ (.CLK(clk),
    .D(_00579_),
    .Q(\data_array.data0[8][37] ));
 sky130_fd_sc_hd__dfxtp_2 _11772_ (.CLK(clk),
    .D(_00580_),
    .Q(\data_array.data0[8][38] ));
 sky130_fd_sc_hd__dfxtp_2 _11773_ (.CLK(clk),
    .D(_00581_),
    .Q(\data_array.data0[8][39] ));
 sky130_fd_sc_hd__dfxtp_2 _11774_ (.CLK(clk),
    .D(_00582_),
    .Q(\data_array.data0[8][40] ));
 sky130_fd_sc_hd__dfxtp_2 _11775_ (.CLK(clk),
    .D(_00583_),
    .Q(\data_array.data0[8][41] ));
 sky130_fd_sc_hd__dfxtp_2 _11776_ (.CLK(clk),
    .D(_00584_),
    .Q(\data_array.data0[8][42] ));
 sky130_fd_sc_hd__dfxtp_2 _11777_ (.CLK(clk),
    .D(_00585_),
    .Q(\data_array.data0[8][43] ));
 sky130_fd_sc_hd__dfxtp_2 _11778_ (.CLK(clk),
    .D(_00586_),
    .Q(\data_array.data0[8][44] ));
 sky130_fd_sc_hd__dfxtp_2 _11779_ (.CLK(clk),
    .D(_00587_),
    .Q(\data_array.data0[8][45] ));
 sky130_fd_sc_hd__dfxtp_2 _11780_ (.CLK(clk),
    .D(_00588_),
    .Q(\data_array.data0[8][46] ));
 sky130_fd_sc_hd__dfxtp_2 _11781_ (.CLK(clk),
    .D(_00589_),
    .Q(\data_array.data0[8][47] ));
 sky130_fd_sc_hd__dfxtp_2 _11782_ (.CLK(clk),
    .D(_00590_),
    .Q(\data_array.data0[8][48] ));
 sky130_fd_sc_hd__dfxtp_2 _11783_ (.CLK(clk),
    .D(_00591_),
    .Q(\data_array.data0[8][49] ));
 sky130_fd_sc_hd__dfxtp_2 _11784_ (.CLK(clk),
    .D(_00592_),
    .Q(\data_array.data0[8][50] ));
 sky130_fd_sc_hd__dfxtp_2 _11785_ (.CLK(clk),
    .D(_00593_),
    .Q(\data_array.data0[8][51] ));
 sky130_fd_sc_hd__dfxtp_2 _11786_ (.CLK(clk),
    .D(_00594_),
    .Q(\data_array.data0[8][52] ));
 sky130_fd_sc_hd__dfxtp_2 _11787_ (.CLK(clk),
    .D(_00595_),
    .Q(\data_array.data0[8][53] ));
 sky130_fd_sc_hd__dfxtp_2 _11788_ (.CLK(clk),
    .D(_00596_),
    .Q(\data_array.data0[8][54] ));
 sky130_fd_sc_hd__dfxtp_2 _11789_ (.CLK(clk),
    .D(_00597_),
    .Q(\data_array.data0[8][55] ));
 sky130_fd_sc_hd__dfxtp_2 _11790_ (.CLK(clk),
    .D(_00598_),
    .Q(\data_array.data0[8][56] ));
 sky130_fd_sc_hd__dfxtp_2 _11791_ (.CLK(clk),
    .D(_00599_),
    .Q(\data_array.data0[8][57] ));
 sky130_fd_sc_hd__dfxtp_2 _11792_ (.CLK(clk),
    .D(_00600_),
    .Q(\data_array.data0[8][58] ));
 sky130_fd_sc_hd__dfxtp_2 _11793_ (.CLK(clk),
    .D(_00601_),
    .Q(\data_array.data0[8][59] ));
 sky130_fd_sc_hd__dfxtp_2 _11794_ (.CLK(clk),
    .D(_00602_),
    .Q(\data_array.data0[8][60] ));
 sky130_fd_sc_hd__dfxtp_2 _11795_ (.CLK(clk),
    .D(_00603_),
    .Q(\data_array.data0[8][61] ));
 sky130_fd_sc_hd__dfxtp_2 _11796_ (.CLK(clk),
    .D(_00604_),
    .Q(\data_array.data0[8][62] ));
 sky130_fd_sc_hd__dfxtp_2 _11797_ (.CLK(clk),
    .D(_00605_),
    .Q(\data_array.data0[8][63] ));
 sky130_fd_sc_hd__dfxtp_2 _11798_ (.CLK(clk),
    .D(_00606_),
    .Q(\data_array.data0[7][0] ));
 sky130_fd_sc_hd__dfxtp_2 _11799_ (.CLK(clk),
    .D(_00607_),
    .Q(\data_array.data0[7][1] ));
 sky130_fd_sc_hd__dfxtp_2 _11800_ (.CLK(clk),
    .D(_00608_),
    .Q(\data_array.data0[7][2] ));
 sky130_fd_sc_hd__dfxtp_2 _11801_ (.CLK(clk),
    .D(_00609_),
    .Q(\data_array.data0[7][3] ));
 sky130_fd_sc_hd__dfxtp_2 _11802_ (.CLK(clk),
    .D(_00610_),
    .Q(\data_array.data0[7][4] ));
 sky130_fd_sc_hd__dfxtp_2 _11803_ (.CLK(clk),
    .D(_00611_),
    .Q(\data_array.data0[7][5] ));
 sky130_fd_sc_hd__dfxtp_2 _11804_ (.CLK(clk),
    .D(_00612_),
    .Q(\data_array.data0[7][6] ));
 sky130_fd_sc_hd__dfxtp_2 _11805_ (.CLK(clk),
    .D(_00613_),
    .Q(\data_array.data0[7][7] ));
 sky130_fd_sc_hd__dfxtp_2 _11806_ (.CLK(clk),
    .D(_00614_),
    .Q(\data_array.data0[7][8] ));
 sky130_fd_sc_hd__dfxtp_2 _11807_ (.CLK(clk),
    .D(_00615_),
    .Q(\data_array.data0[7][9] ));
 sky130_fd_sc_hd__dfxtp_2 _11808_ (.CLK(clk),
    .D(_00616_),
    .Q(\data_array.data0[7][10] ));
 sky130_fd_sc_hd__dfxtp_2 _11809_ (.CLK(clk),
    .D(_00617_),
    .Q(\data_array.data0[7][11] ));
 sky130_fd_sc_hd__dfxtp_2 _11810_ (.CLK(clk),
    .D(_00618_),
    .Q(\data_array.data0[7][12] ));
 sky130_fd_sc_hd__dfxtp_2 _11811_ (.CLK(clk),
    .D(_00619_),
    .Q(\data_array.data0[7][13] ));
 sky130_fd_sc_hd__dfxtp_2 _11812_ (.CLK(clk),
    .D(_00620_),
    .Q(\data_array.data0[7][14] ));
 sky130_fd_sc_hd__dfxtp_2 _11813_ (.CLK(clk),
    .D(_00621_),
    .Q(\data_array.data0[7][15] ));
 sky130_fd_sc_hd__dfxtp_2 _11814_ (.CLK(clk),
    .D(_00622_),
    .Q(\data_array.data0[7][16] ));
 sky130_fd_sc_hd__dfxtp_2 _11815_ (.CLK(clk),
    .D(_00623_),
    .Q(\data_array.data0[7][17] ));
 sky130_fd_sc_hd__dfxtp_2 _11816_ (.CLK(clk),
    .D(_00624_),
    .Q(\data_array.data0[7][18] ));
 sky130_fd_sc_hd__dfxtp_2 _11817_ (.CLK(clk),
    .D(_00625_),
    .Q(\data_array.data0[7][19] ));
 sky130_fd_sc_hd__dfxtp_2 _11818_ (.CLK(clk),
    .D(_00626_),
    .Q(\data_array.data0[7][20] ));
 sky130_fd_sc_hd__dfxtp_2 _11819_ (.CLK(clk),
    .D(_00627_),
    .Q(\data_array.data0[7][21] ));
 sky130_fd_sc_hd__dfxtp_2 _11820_ (.CLK(clk),
    .D(_00628_),
    .Q(\data_array.data0[7][22] ));
 sky130_fd_sc_hd__dfxtp_2 _11821_ (.CLK(clk),
    .D(_00629_),
    .Q(\data_array.data0[7][23] ));
 sky130_fd_sc_hd__dfxtp_2 _11822_ (.CLK(clk),
    .D(_00630_),
    .Q(\data_array.data0[7][24] ));
 sky130_fd_sc_hd__dfxtp_2 _11823_ (.CLK(clk),
    .D(_00631_),
    .Q(\data_array.data0[7][25] ));
 sky130_fd_sc_hd__dfxtp_2 _11824_ (.CLK(clk),
    .D(_00632_),
    .Q(\data_array.data0[7][26] ));
 sky130_fd_sc_hd__dfxtp_2 _11825_ (.CLK(clk),
    .D(_00633_),
    .Q(\data_array.data0[7][27] ));
 sky130_fd_sc_hd__dfxtp_2 _11826_ (.CLK(clk),
    .D(_00634_),
    .Q(\data_array.data0[7][28] ));
 sky130_fd_sc_hd__dfxtp_2 _11827_ (.CLK(clk),
    .D(_00635_),
    .Q(\data_array.data0[7][29] ));
 sky130_fd_sc_hd__dfxtp_2 _11828_ (.CLK(clk),
    .D(_00636_),
    .Q(\data_array.data0[7][30] ));
 sky130_fd_sc_hd__dfxtp_2 _11829_ (.CLK(clk),
    .D(_00637_),
    .Q(\data_array.data0[7][31] ));
 sky130_fd_sc_hd__dfxtp_2 _11830_ (.CLK(clk),
    .D(_00638_),
    .Q(\data_array.data0[7][32] ));
 sky130_fd_sc_hd__dfxtp_2 _11831_ (.CLK(clk),
    .D(_00639_),
    .Q(\data_array.data0[7][33] ));
 sky130_fd_sc_hd__dfxtp_2 _11832_ (.CLK(clk),
    .D(_00640_),
    .Q(\data_array.data0[7][34] ));
 sky130_fd_sc_hd__dfxtp_2 _11833_ (.CLK(clk),
    .D(_00641_),
    .Q(\data_array.data0[7][35] ));
 sky130_fd_sc_hd__dfxtp_2 _11834_ (.CLK(clk),
    .D(_00642_),
    .Q(\data_array.data0[7][36] ));
 sky130_fd_sc_hd__dfxtp_2 _11835_ (.CLK(clk),
    .D(_00643_),
    .Q(\data_array.data0[7][37] ));
 sky130_fd_sc_hd__dfxtp_2 _11836_ (.CLK(clk),
    .D(_00644_),
    .Q(\data_array.data0[7][38] ));
 sky130_fd_sc_hd__dfxtp_2 _11837_ (.CLK(clk),
    .D(_00645_),
    .Q(\data_array.data0[7][39] ));
 sky130_fd_sc_hd__dfxtp_2 _11838_ (.CLK(clk),
    .D(_00646_),
    .Q(\data_array.data0[7][40] ));
 sky130_fd_sc_hd__dfxtp_2 _11839_ (.CLK(clk),
    .D(_00647_),
    .Q(\data_array.data0[7][41] ));
 sky130_fd_sc_hd__dfxtp_2 _11840_ (.CLK(clk),
    .D(_00648_),
    .Q(\data_array.data0[7][42] ));
 sky130_fd_sc_hd__dfxtp_2 _11841_ (.CLK(clk),
    .D(_00649_),
    .Q(\data_array.data0[7][43] ));
 sky130_fd_sc_hd__dfxtp_2 _11842_ (.CLK(clk),
    .D(_00650_),
    .Q(\data_array.data0[7][44] ));
 sky130_fd_sc_hd__dfxtp_2 _11843_ (.CLK(clk),
    .D(_00651_),
    .Q(\data_array.data0[7][45] ));
 sky130_fd_sc_hd__dfxtp_2 _11844_ (.CLK(clk),
    .D(_00652_),
    .Q(\data_array.data0[7][46] ));
 sky130_fd_sc_hd__dfxtp_2 _11845_ (.CLK(clk),
    .D(_00653_),
    .Q(\data_array.data0[7][47] ));
 sky130_fd_sc_hd__dfxtp_2 _11846_ (.CLK(clk),
    .D(_00654_),
    .Q(\data_array.data0[7][48] ));
 sky130_fd_sc_hd__dfxtp_2 _11847_ (.CLK(clk),
    .D(_00655_),
    .Q(\data_array.data0[7][49] ));
 sky130_fd_sc_hd__dfxtp_2 _11848_ (.CLK(clk),
    .D(_00656_),
    .Q(\data_array.data0[7][50] ));
 sky130_fd_sc_hd__dfxtp_2 _11849_ (.CLK(clk),
    .D(_00657_),
    .Q(\data_array.data0[7][51] ));
 sky130_fd_sc_hd__dfxtp_2 _11850_ (.CLK(clk),
    .D(_00658_),
    .Q(\data_array.data0[7][52] ));
 sky130_fd_sc_hd__dfxtp_2 _11851_ (.CLK(clk),
    .D(_00659_),
    .Q(\data_array.data0[7][53] ));
 sky130_fd_sc_hd__dfxtp_2 _11852_ (.CLK(clk),
    .D(_00660_),
    .Q(\data_array.data0[7][54] ));
 sky130_fd_sc_hd__dfxtp_2 _11853_ (.CLK(clk),
    .D(_00661_),
    .Q(\data_array.data0[7][55] ));
 sky130_fd_sc_hd__dfxtp_2 _11854_ (.CLK(clk),
    .D(_00662_),
    .Q(\data_array.data0[7][56] ));
 sky130_fd_sc_hd__dfxtp_2 _11855_ (.CLK(clk),
    .D(_00663_),
    .Q(\data_array.data0[7][57] ));
 sky130_fd_sc_hd__dfxtp_2 _11856_ (.CLK(clk),
    .D(_00664_),
    .Q(\data_array.data0[7][58] ));
 sky130_fd_sc_hd__dfxtp_2 _11857_ (.CLK(clk),
    .D(_00665_),
    .Q(\data_array.data0[7][59] ));
 sky130_fd_sc_hd__dfxtp_2 _11858_ (.CLK(clk),
    .D(_00666_),
    .Q(\data_array.data0[7][60] ));
 sky130_fd_sc_hd__dfxtp_2 _11859_ (.CLK(clk),
    .D(_00667_),
    .Q(\data_array.data0[7][61] ));
 sky130_fd_sc_hd__dfxtp_2 _11860_ (.CLK(clk),
    .D(_00668_),
    .Q(\data_array.data0[7][62] ));
 sky130_fd_sc_hd__dfxtp_2 _11861_ (.CLK(clk),
    .D(_00669_),
    .Q(\data_array.data0[7][63] ));
 sky130_fd_sc_hd__dfxtp_2 _11862_ (.CLK(clk),
    .D(_00670_),
    .Q(\data_array.data0[5][0] ));
 sky130_fd_sc_hd__dfxtp_2 _11863_ (.CLK(clk),
    .D(_00671_),
    .Q(\data_array.data0[5][1] ));
 sky130_fd_sc_hd__dfxtp_2 _11864_ (.CLK(clk),
    .D(_00672_),
    .Q(\data_array.data0[5][2] ));
 sky130_fd_sc_hd__dfxtp_2 _11865_ (.CLK(clk),
    .D(_00673_),
    .Q(\data_array.data0[5][3] ));
 sky130_fd_sc_hd__dfxtp_2 _11866_ (.CLK(clk),
    .D(_00674_),
    .Q(\data_array.data0[5][4] ));
 sky130_fd_sc_hd__dfxtp_2 _11867_ (.CLK(clk),
    .D(_00675_),
    .Q(\data_array.data0[5][5] ));
 sky130_fd_sc_hd__dfxtp_2 _11868_ (.CLK(clk),
    .D(_00676_),
    .Q(\data_array.data0[5][6] ));
 sky130_fd_sc_hd__dfxtp_2 _11869_ (.CLK(clk),
    .D(_00677_),
    .Q(\data_array.data0[5][7] ));
 sky130_fd_sc_hd__dfxtp_2 _11870_ (.CLK(clk),
    .D(_00678_),
    .Q(\data_array.data0[5][8] ));
 sky130_fd_sc_hd__dfxtp_2 _11871_ (.CLK(clk),
    .D(_00679_),
    .Q(\data_array.data0[5][9] ));
 sky130_fd_sc_hd__dfxtp_2 _11872_ (.CLK(clk),
    .D(_00680_),
    .Q(\data_array.data0[5][10] ));
 sky130_fd_sc_hd__dfxtp_2 _11873_ (.CLK(clk),
    .D(_00681_),
    .Q(\data_array.data0[5][11] ));
 sky130_fd_sc_hd__dfxtp_2 _11874_ (.CLK(clk),
    .D(_00682_),
    .Q(\data_array.data0[5][12] ));
 sky130_fd_sc_hd__dfxtp_2 _11875_ (.CLK(clk),
    .D(_00683_),
    .Q(\data_array.data0[5][13] ));
 sky130_fd_sc_hd__dfxtp_2 _11876_ (.CLK(clk),
    .D(_00684_),
    .Q(\data_array.data0[5][14] ));
 sky130_fd_sc_hd__dfxtp_2 _11877_ (.CLK(clk),
    .D(_00685_),
    .Q(\data_array.data0[5][15] ));
 sky130_fd_sc_hd__dfxtp_2 _11878_ (.CLK(clk),
    .D(_00686_),
    .Q(\data_array.data0[5][16] ));
 sky130_fd_sc_hd__dfxtp_2 _11879_ (.CLK(clk),
    .D(_00687_),
    .Q(\data_array.data0[5][17] ));
 sky130_fd_sc_hd__dfxtp_2 _11880_ (.CLK(clk),
    .D(_00688_),
    .Q(\data_array.data0[5][18] ));
 sky130_fd_sc_hd__dfxtp_2 _11881_ (.CLK(clk),
    .D(_00689_),
    .Q(\data_array.data0[5][19] ));
 sky130_fd_sc_hd__dfxtp_2 _11882_ (.CLK(clk),
    .D(_00690_),
    .Q(\data_array.data0[5][20] ));
 sky130_fd_sc_hd__dfxtp_2 _11883_ (.CLK(clk),
    .D(_00691_),
    .Q(\data_array.data0[5][21] ));
 sky130_fd_sc_hd__dfxtp_2 _11884_ (.CLK(clk),
    .D(_00692_),
    .Q(\data_array.data0[5][22] ));
 sky130_fd_sc_hd__dfxtp_2 _11885_ (.CLK(clk),
    .D(_00693_),
    .Q(\data_array.data0[5][23] ));
 sky130_fd_sc_hd__dfxtp_2 _11886_ (.CLK(clk),
    .D(_00694_),
    .Q(\data_array.data0[5][24] ));
 sky130_fd_sc_hd__dfxtp_2 _11887_ (.CLK(clk),
    .D(_00695_),
    .Q(\data_array.data0[5][25] ));
 sky130_fd_sc_hd__dfxtp_2 _11888_ (.CLK(clk),
    .D(_00696_),
    .Q(\data_array.data0[5][26] ));
 sky130_fd_sc_hd__dfxtp_2 _11889_ (.CLK(clk),
    .D(_00697_),
    .Q(\data_array.data0[5][27] ));
 sky130_fd_sc_hd__dfxtp_2 _11890_ (.CLK(clk),
    .D(_00698_),
    .Q(\data_array.data0[5][28] ));
 sky130_fd_sc_hd__dfxtp_2 _11891_ (.CLK(clk),
    .D(_00699_),
    .Q(\data_array.data0[5][29] ));
 sky130_fd_sc_hd__dfxtp_2 _11892_ (.CLK(clk),
    .D(_00700_),
    .Q(\data_array.data0[5][30] ));
 sky130_fd_sc_hd__dfxtp_2 _11893_ (.CLK(clk),
    .D(_00701_),
    .Q(\data_array.data0[5][31] ));
 sky130_fd_sc_hd__dfxtp_2 _11894_ (.CLK(clk),
    .D(_00702_),
    .Q(\data_array.data0[5][32] ));
 sky130_fd_sc_hd__dfxtp_2 _11895_ (.CLK(clk),
    .D(_00703_),
    .Q(\data_array.data0[5][33] ));
 sky130_fd_sc_hd__dfxtp_2 _11896_ (.CLK(clk),
    .D(_00704_),
    .Q(\data_array.data0[5][34] ));
 sky130_fd_sc_hd__dfxtp_2 _11897_ (.CLK(clk),
    .D(_00705_),
    .Q(\data_array.data0[5][35] ));
 sky130_fd_sc_hd__dfxtp_2 _11898_ (.CLK(clk),
    .D(_00706_),
    .Q(\data_array.data0[5][36] ));
 sky130_fd_sc_hd__dfxtp_2 _11899_ (.CLK(clk),
    .D(_00707_),
    .Q(\data_array.data0[5][37] ));
 sky130_fd_sc_hd__dfxtp_2 _11900_ (.CLK(clk),
    .D(_00708_),
    .Q(\data_array.data0[5][38] ));
 sky130_fd_sc_hd__dfxtp_2 _11901_ (.CLK(clk),
    .D(_00709_),
    .Q(\data_array.data0[5][39] ));
 sky130_fd_sc_hd__dfxtp_2 _11902_ (.CLK(clk),
    .D(_00710_),
    .Q(\data_array.data0[5][40] ));
 sky130_fd_sc_hd__dfxtp_2 _11903_ (.CLK(clk),
    .D(_00711_),
    .Q(\data_array.data0[5][41] ));
 sky130_fd_sc_hd__dfxtp_2 _11904_ (.CLK(clk),
    .D(_00712_),
    .Q(\data_array.data0[5][42] ));
 sky130_fd_sc_hd__dfxtp_2 _11905_ (.CLK(clk),
    .D(_00713_),
    .Q(\data_array.data0[5][43] ));
 sky130_fd_sc_hd__dfxtp_2 _11906_ (.CLK(clk),
    .D(_00714_),
    .Q(\data_array.data0[5][44] ));
 sky130_fd_sc_hd__dfxtp_2 _11907_ (.CLK(clk),
    .D(_00715_),
    .Q(\data_array.data0[5][45] ));
 sky130_fd_sc_hd__dfxtp_2 _11908_ (.CLK(clk),
    .D(_00716_),
    .Q(\data_array.data0[5][46] ));
 sky130_fd_sc_hd__dfxtp_2 _11909_ (.CLK(clk),
    .D(_00717_),
    .Q(\data_array.data0[5][47] ));
 sky130_fd_sc_hd__dfxtp_2 _11910_ (.CLK(clk),
    .D(_00718_),
    .Q(\data_array.data0[5][48] ));
 sky130_fd_sc_hd__dfxtp_2 _11911_ (.CLK(clk),
    .D(_00719_),
    .Q(\data_array.data0[5][49] ));
 sky130_fd_sc_hd__dfxtp_2 _11912_ (.CLK(clk),
    .D(_00720_),
    .Q(\data_array.data0[5][50] ));
 sky130_fd_sc_hd__dfxtp_2 _11913_ (.CLK(clk),
    .D(_00721_),
    .Q(\data_array.data0[5][51] ));
 sky130_fd_sc_hd__dfxtp_2 _11914_ (.CLK(clk),
    .D(_00722_),
    .Q(\data_array.data0[5][52] ));
 sky130_fd_sc_hd__dfxtp_2 _11915_ (.CLK(clk),
    .D(_00723_),
    .Q(\data_array.data0[5][53] ));
 sky130_fd_sc_hd__dfxtp_2 _11916_ (.CLK(clk),
    .D(_00724_),
    .Q(\data_array.data0[5][54] ));
 sky130_fd_sc_hd__dfxtp_2 _11917_ (.CLK(clk),
    .D(_00725_),
    .Q(\data_array.data0[5][55] ));
 sky130_fd_sc_hd__dfxtp_2 _11918_ (.CLK(clk),
    .D(_00726_),
    .Q(\data_array.data0[5][56] ));
 sky130_fd_sc_hd__dfxtp_2 _11919_ (.CLK(clk),
    .D(_00727_),
    .Q(\data_array.data0[5][57] ));
 sky130_fd_sc_hd__dfxtp_2 _11920_ (.CLK(clk),
    .D(_00728_),
    .Q(\data_array.data0[5][58] ));
 sky130_fd_sc_hd__dfxtp_2 _11921_ (.CLK(clk),
    .D(_00729_),
    .Q(\data_array.data0[5][59] ));
 sky130_fd_sc_hd__dfxtp_2 _11922_ (.CLK(clk),
    .D(_00730_),
    .Q(\data_array.data0[5][60] ));
 sky130_fd_sc_hd__dfxtp_2 _11923_ (.CLK(clk),
    .D(_00731_),
    .Q(\data_array.data0[5][61] ));
 sky130_fd_sc_hd__dfxtp_2 _11924_ (.CLK(clk),
    .D(_00732_),
    .Q(\data_array.data0[5][62] ));
 sky130_fd_sc_hd__dfxtp_2 _11925_ (.CLK(clk),
    .D(_00733_),
    .Q(\data_array.data0[5][63] ));
 sky130_fd_sc_hd__dfxtp_2 _11926_ (.CLK(clk),
    .D(_00734_),
    .Q(\data_array.data0[4][0] ));
 sky130_fd_sc_hd__dfxtp_2 _11927_ (.CLK(clk),
    .D(_00735_),
    .Q(\data_array.data0[4][1] ));
 sky130_fd_sc_hd__dfxtp_2 _11928_ (.CLK(clk),
    .D(_00736_),
    .Q(\data_array.data0[4][2] ));
 sky130_fd_sc_hd__dfxtp_2 _11929_ (.CLK(clk),
    .D(_00737_),
    .Q(\data_array.data0[4][3] ));
 sky130_fd_sc_hd__dfxtp_2 _11930_ (.CLK(clk),
    .D(_00738_),
    .Q(\data_array.data0[4][4] ));
 sky130_fd_sc_hd__dfxtp_2 _11931_ (.CLK(clk),
    .D(_00739_),
    .Q(\data_array.data0[4][5] ));
 sky130_fd_sc_hd__dfxtp_2 _11932_ (.CLK(clk),
    .D(_00740_),
    .Q(\data_array.data0[4][6] ));
 sky130_fd_sc_hd__dfxtp_2 _11933_ (.CLK(clk),
    .D(_00741_),
    .Q(\data_array.data0[4][7] ));
 sky130_fd_sc_hd__dfxtp_2 _11934_ (.CLK(clk),
    .D(_00742_),
    .Q(\data_array.data0[4][8] ));
 sky130_fd_sc_hd__dfxtp_2 _11935_ (.CLK(clk),
    .D(_00743_),
    .Q(\data_array.data0[4][9] ));
 sky130_fd_sc_hd__dfxtp_2 _11936_ (.CLK(clk),
    .D(_00744_),
    .Q(\data_array.data0[4][10] ));
 sky130_fd_sc_hd__dfxtp_2 _11937_ (.CLK(clk),
    .D(_00745_),
    .Q(\data_array.data0[4][11] ));
 sky130_fd_sc_hd__dfxtp_2 _11938_ (.CLK(clk),
    .D(_00746_),
    .Q(\data_array.data0[4][12] ));
 sky130_fd_sc_hd__dfxtp_2 _11939_ (.CLK(clk),
    .D(_00747_),
    .Q(\data_array.data0[4][13] ));
 sky130_fd_sc_hd__dfxtp_2 _11940_ (.CLK(clk),
    .D(_00748_),
    .Q(\data_array.data0[4][14] ));
 sky130_fd_sc_hd__dfxtp_2 _11941_ (.CLK(clk),
    .D(_00749_),
    .Q(\data_array.data0[4][15] ));
 sky130_fd_sc_hd__dfxtp_2 _11942_ (.CLK(clk),
    .D(_00750_),
    .Q(\data_array.data0[4][16] ));
 sky130_fd_sc_hd__dfxtp_2 _11943_ (.CLK(clk),
    .D(_00751_),
    .Q(\data_array.data0[4][17] ));
 sky130_fd_sc_hd__dfxtp_2 _11944_ (.CLK(clk),
    .D(_00752_),
    .Q(\data_array.data0[4][18] ));
 sky130_fd_sc_hd__dfxtp_2 _11945_ (.CLK(clk),
    .D(_00753_),
    .Q(\data_array.data0[4][19] ));
 sky130_fd_sc_hd__dfxtp_2 _11946_ (.CLK(clk),
    .D(_00754_),
    .Q(\data_array.data0[4][20] ));
 sky130_fd_sc_hd__dfxtp_2 _11947_ (.CLK(clk),
    .D(_00755_),
    .Q(\data_array.data0[4][21] ));
 sky130_fd_sc_hd__dfxtp_2 _11948_ (.CLK(clk),
    .D(_00756_),
    .Q(\data_array.data0[4][22] ));
 sky130_fd_sc_hd__dfxtp_2 _11949_ (.CLK(clk),
    .D(_00757_),
    .Q(\data_array.data0[4][23] ));
 sky130_fd_sc_hd__dfxtp_2 _11950_ (.CLK(clk),
    .D(_00758_),
    .Q(\data_array.data0[4][24] ));
 sky130_fd_sc_hd__dfxtp_2 _11951_ (.CLK(clk),
    .D(_00759_),
    .Q(\data_array.data0[4][25] ));
 sky130_fd_sc_hd__dfxtp_2 _11952_ (.CLK(clk),
    .D(_00760_),
    .Q(\data_array.data0[4][26] ));
 sky130_fd_sc_hd__dfxtp_2 _11953_ (.CLK(clk),
    .D(_00761_),
    .Q(\data_array.data0[4][27] ));
 sky130_fd_sc_hd__dfxtp_2 _11954_ (.CLK(clk),
    .D(_00762_),
    .Q(\data_array.data0[4][28] ));
 sky130_fd_sc_hd__dfxtp_2 _11955_ (.CLK(clk),
    .D(_00763_),
    .Q(\data_array.data0[4][29] ));
 sky130_fd_sc_hd__dfxtp_2 _11956_ (.CLK(clk),
    .D(_00764_),
    .Q(\data_array.data0[4][30] ));
 sky130_fd_sc_hd__dfxtp_2 _11957_ (.CLK(clk),
    .D(_00765_),
    .Q(\data_array.data0[4][31] ));
 sky130_fd_sc_hd__dfxtp_2 _11958_ (.CLK(clk),
    .D(_00766_),
    .Q(\data_array.data0[4][32] ));
 sky130_fd_sc_hd__dfxtp_2 _11959_ (.CLK(clk),
    .D(_00767_),
    .Q(\data_array.data0[4][33] ));
 sky130_fd_sc_hd__dfxtp_2 _11960_ (.CLK(clk),
    .D(_00768_),
    .Q(\data_array.data0[4][34] ));
 sky130_fd_sc_hd__dfxtp_2 _11961_ (.CLK(clk),
    .D(_00769_),
    .Q(\data_array.data0[4][35] ));
 sky130_fd_sc_hd__dfxtp_2 _11962_ (.CLK(clk),
    .D(_00770_),
    .Q(\data_array.data0[4][36] ));
 sky130_fd_sc_hd__dfxtp_2 _11963_ (.CLK(clk),
    .D(_00771_),
    .Q(\data_array.data0[4][37] ));
 sky130_fd_sc_hd__dfxtp_2 _11964_ (.CLK(clk),
    .D(_00772_),
    .Q(\data_array.data0[4][38] ));
 sky130_fd_sc_hd__dfxtp_2 _11965_ (.CLK(clk),
    .D(_00773_),
    .Q(\data_array.data0[4][39] ));
 sky130_fd_sc_hd__dfxtp_2 _11966_ (.CLK(clk),
    .D(_00774_),
    .Q(\data_array.data0[4][40] ));
 sky130_fd_sc_hd__dfxtp_2 _11967_ (.CLK(clk),
    .D(_00775_),
    .Q(\data_array.data0[4][41] ));
 sky130_fd_sc_hd__dfxtp_2 _11968_ (.CLK(clk),
    .D(_00776_),
    .Q(\data_array.data0[4][42] ));
 sky130_fd_sc_hd__dfxtp_2 _11969_ (.CLK(clk),
    .D(_00777_),
    .Q(\data_array.data0[4][43] ));
 sky130_fd_sc_hd__dfxtp_2 _11970_ (.CLK(clk),
    .D(_00778_),
    .Q(\data_array.data0[4][44] ));
 sky130_fd_sc_hd__dfxtp_2 _11971_ (.CLK(clk),
    .D(_00779_),
    .Q(\data_array.data0[4][45] ));
 sky130_fd_sc_hd__dfxtp_2 _11972_ (.CLK(clk),
    .D(_00780_),
    .Q(\data_array.data0[4][46] ));
 sky130_fd_sc_hd__dfxtp_2 _11973_ (.CLK(clk),
    .D(_00781_),
    .Q(\data_array.data0[4][47] ));
 sky130_fd_sc_hd__dfxtp_2 _11974_ (.CLK(clk),
    .D(_00782_),
    .Q(\data_array.data0[4][48] ));
 sky130_fd_sc_hd__dfxtp_2 _11975_ (.CLK(clk),
    .D(_00783_),
    .Q(\data_array.data0[4][49] ));
 sky130_fd_sc_hd__dfxtp_2 _11976_ (.CLK(clk),
    .D(_00784_),
    .Q(\data_array.data0[4][50] ));
 sky130_fd_sc_hd__dfxtp_2 _11977_ (.CLK(clk),
    .D(_00785_),
    .Q(\data_array.data0[4][51] ));
 sky130_fd_sc_hd__dfxtp_2 _11978_ (.CLK(clk),
    .D(_00786_),
    .Q(\data_array.data0[4][52] ));
 sky130_fd_sc_hd__dfxtp_2 _11979_ (.CLK(clk),
    .D(_00787_),
    .Q(\data_array.data0[4][53] ));
 sky130_fd_sc_hd__dfxtp_2 _11980_ (.CLK(clk),
    .D(_00788_),
    .Q(\data_array.data0[4][54] ));
 sky130_fd_sc_hd__dfxtp_2 _11981_ (.CLK(clk),
    .D(_00789_),
    .Q(\data_array.data0[4][55] ));
 sky130_fd_sc_hd__dfxtp_2 _11982_ (.CLK(clk),
    .D(_00790_),
    .Q(\data_array.data0[4][56] ));
 sky130_fd_sc_hd__dfxtp_2 _11983_ (.CLK(clk),
    .D(_00791_),
    .Q(\data_array.data0[4][57] ));
 sky130_fd_sc_hd__dfxtp_2 _11984_ (.CLK(clk),
    .D(_00792_),
    .Q(\data_array.data0[4][58] ));
 sky130_fd_sc_hd__dfxtp_2 _11985_ (.CLK(clk),
    .D(_00793_),
    .Q(\data_array.data0[4][59] ));
 sky130_fd_sc_hd__dfxtp_2 _11986_ (.CLK(clk),
    .D(_00794_),
    .Q(\data_array.data0[4][60] ));
 sky130_fd_sc_hd__dfxtp_2 _11987_ (.CLK(clk),
    .D(_00795_),
    .Q(\data_array.data0[4][61] ));
 sky130_fd_sc_hd__dfxtp_2 _11988_ (.CLK(clk),
    .D(_00796_),
    .Q(\data_array.data0[4][62] ));
 sky130_fd_sc_hd__dfxtp_2 _11989_ (.CLK(clk),
    .D(_00797_),
    .Q(\data_array.data0[4][63] ));
 sky130_fd_sc_hd__dfxtp_2 _11990_ (.CLK(clk),
    .D(_00798_),
    .Q(\data_array.data0[6][0] ));
 sky130_fd_sc_hd__dfxtp_2 _11991_ (.CLK(clk),
    .D(_00799_),
    .Q(\data_array.data0[6][1] ));
 sky130_fd_sc_hd__dfxtp_2 _11992_ (.CLK(clk),
    .D(_00800_),
    .Q(\data_array.data0[6][2] ));
 sky130_fd_sc_hd__dfxtp_2 _11993_ (.CLK(clk),
    .D(_00801_),
    .Q(\data_array.data0[6][3] ));
 sky130_fd_sc_hd__dfxtp_2 _11994_ (.CLK(clk),
    .D(_00802_),
    .Q(\data_array.data0[6][4] ));
 sky130_fd_sc_hd__dfxtp_2 _11995_ (.CLK(clk),
    .D(_00803_),
    .Q(\data_array.data0[6][5] ));
 sky130_fd_sc_hd__dfxtp_2 _11996_ (.CLK(clk),
    .D(_00804_),
    .Q(\data_array.data0[6][6] ));
 sky130_fd_sc_hd__dfxtp_2 _11997_ (.CLK(clk),
    .D(_00805_),
    .Q(\data_array.data0[6][7] ));
 sky130_fd_sc_hd__dfxtp_2 _11998_ (.CLK(clk),
    .D(_00806_),
    .Q(\data_array.data0[6][8] ));
 sky130_fd_sc_hd__dfxtp_2 _11999_ (.CLK(clk),
    .D(_00807_),
    .Q(\data_array.data0[6][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12000_ (.CLK(clk),
    .D(_00808_),
    .Q(\data_array.data0[6][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12001_ (.CLK(clk),
    .D(_00809_),
    .Q(\data_array.data0[6][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12002_ (.CLK(clk),
    .D(_00810_),
    .Q(\data_array.data0[6][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12003_ (.CLK(clk),
    .D(_00811_),
    .Q(\data_array.data0[6][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12004_ (.CLK(clk),
    .D(_00812_),
    .Q(\data_array.data0[6][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12005_ (.CLK(clk),
    .D(_00813_),
    .Q(\data_array.data0[6][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12006_ (.CLK(clk),
    .D(_00814_),
    .Q(\data_array.data0[6][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12007_ (.CLK(clk),
    .D(_00815_),
    .Q(\data_array.data0[6][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12008_ (.CLK(clk),
    .D(_00816_),
    .Q(\data_array.data0[6][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12009_ (.CLK(clk),
    .D(_00817_),
    .Q(\data_array.data0[6][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12010_ (.CLK(clk),
    .D(_00818_),
    .Q(\data_array.data0[6][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12011_ (.CLK(clk),
    .D(_00819_),
    .Q(\data_array.data0[6][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12012_ (.CLK(clk),
    .D(_00820_),
    .Q(\data_array.data0[6][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12013_ (.CLK(clk),
    .D(_00821_),
    .Q(\data_array.data0[6][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12014_ (.CLK(clk),
    .D(_00822_),
    .Q(\data_array.data0[6][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12015_ (.CLK(clk),
    .D(_00823_),
    .Q(\data_array.data0[6][25] ));
 sky130_fd_sc_hd__dfxtp_2 _12016_ (.CLK(clk),
    .D(_00824_),
    .Q(\data_array.data0[6][26] ));
 sky130_fd_sc_hd__dfxtp_2 _12017_ (.CLK(clk),
    .D(_00825_),
    .Q(\data_array.data0[6][27] ));
 sky130_fd_sc_hd__dfxtp_2 _12018_ (.CLK(clk),
    .D(_00826_),
    .Q(\data_array.data0[6][28] ));
 sky130_fd_sc_hd__dfxtp_2 _12019_ (.CLK(clk),
    .D(_00827_),
    .Q(\data_array.data0[6][29] ));
 sky130_fd_sc_hd__dfxtp_2 _12020_ (.CLK(clk),
    .D(_00828_),
    .Q(\data_array.data0[6][30] ));
 sky130_fd_sc_hd__dfxtp_2 _12021_ (.CLK(clk),
    .D(_00829_),
    .Q(\data_array.data0[6][31] ));
 sky130_fd_sc_hd__dfxtp_2 _12022_ (.CLK(clk),
    .D(_00830_),
    .Q(\data_array.data0[6][32] ));
 sky130_fd_sc_hd__dfxtp_2 _12023_ (.CLK(clk),
    .D(_00831_),
    .Q(\data_array.data0[6][33] ));
 sky130_fd_sc_hd__dfxtp_2 _12024_ (.CLK(clk),
    .D(_00832_),
    .Q(\data_array.data0[6][34] ));
 sky130_fd_sc_hd__dfxtp_2 _12025_ (.CLK(clk),
    .D(_00833_),
    .Q(\data_array.data0[6][35] ));
 sky130_fd_sc_hd__dfxtp_2 _12026_ (.CLK(clk),
    .D(_00834_),
    .Q(\data_array.data0[6][36] ));
 sky130_fd_sc_hd__dfxtp_2 _12027_ (.CLK(clk),
    .D(_00835_),
    .Q(\data_array.data0[6][37] ));
 sky130_fd_sc_hd__dfxtp_2 _12028_ (.CLK(clk),
    .D(_00836_),
    .Q(\data_array.data0[6][38] ));
 sky130_fd_sc_hd__dfxtp_2 _12029_ (.CLK(clk),
    .D(_00837_),
    .Q(\data_array.data0[6][39] ));
 sky130_fd_sc_hd__dfxtp_2 _12030_ (.CLK(clk),
    .D(_00838_),
    .Q(\data_array.data0[6][40] ));
 sky130_fd_sc_hd__dfxtp_2 _12031_ (.CLK(clk),
    .D(_00839_),
    .Q(\data_array.data0[6][41] ));
 sky130_fd_sc_hd__dfxtp_2 _12032_ (.CLK(clk),
    .D(_00840_),
    .Q(\data_array.data0[6][42] ));
 sky130_fd_sc_hd__dfxtp_2 _12033_ (.CLK(clk),
    .D(_00841_),
    .Q(\data_array.data0[6][43] ));
 sky130_fd_sc_hd__dfxtp_2 _12034_ (.CLK(clk),
    .D(_00842_),
    .Q(\data_array.data0[6][44] ));
 sky130_fd_sc_hd__dfxtp_2 _12035_ (.CLK(clk),
    .D(_00843_),
    .Q(\data_array.data0[6][45] ));
 sky130_fd_sc_hd__dfxtp_2 _12036_ (.CLK(clk),
    .D(_00844_),
    .Q(\data_array.data0[6][46] ));
 sky130_fd_sc_hd__dfxtp_2 _12037_ (.CLK(clk),
    .D(_00845_),
    .Q(\data_array.data0[6][47] ));
 sky130_fd_sc_hd__dfxtp_2 _12038_ (.CLK(clk),
    .D(_00846_),
    .Q(\data_array.data0[6][48] ));
 sky130_fd_sc_hd__dfxtp_2 _12039_ (.CLK(clk),
    .D(_00847_),
    .Q(\data_array.data0[6][49] ));
 sky130_fd_sc_hd__dfxtp_2 _12040_ (.CLK(clk),
    .D(_00848_),
    .Q(\data_array.data0[6][50] ));
 sky130_fd_sc_hd__dfxtp_2 _12041_ (.CLK(clk),
    .D(_00849_),
    .Q(\data_array.data0[6][51] ));
 sky130_fd_sc_hd__dfxtp_2 _12042_ (.CLK(clk),
    .D(_00850_),
    .Q(\data_array.data0[6][52] ));
 sky130_fd_sc_hd__dfxtp_2 _12043_ (.CLK(clk),
    .D(_00851_),
    .Q(\data_array.data0[6][53] ));
 sky130_fd_sc_hd__dfxtp_2 _12044_ (.CLK(clk),
    .D(_00852_),
    .Q(\data_array.data0[6][54] ));
 sky130_fd_sc_hd__dfxtp_2 _12045_ (.CLK(clk),
    .D(_00853_),
    .Q(\data_array.data0[6][55] ));
 sky130_fd_sc_hd__dfxtp_2 _12046_ (.CLK(clk),
    .D(_00854_),
    .Q(\data_array.data0[6][56] ));
 sky130_fd_sc_hd__dfxtp_2 _12047_ (.CLK(clk),
    .D(_00855_),
    .Q(\data_array.data0[6][57] ));
 sky130_fd_sc_hd__dfxtp_2 _12048_ (.CLK(clk),
    .D(_00856_),
    .Q(\data_array.data0[6][58] ));
 sky130_fd_sc_hd__dfxtp_2 _12049_ (.CLK(clk),
    .D(_00857_),
    .Q(\data_array.data0[6][59] ));
 sky130_fd_sc_hd__dfxtp_2 _12050_ (.CLK(clk),
    .D(_00858_),
    .Q(\data_array.data0[6][60] ));
 sky130_fd_sc_hd__dfxtp_2 _12051_ (.CLK(clk),
    .D(_00859_),
    .Q(\data_array.data0[6][61] ));
 sky130_fd_sc_hd__dfxtp_2 _12052_ (.CLK(clk),
    .D(_00860_),
    .Q(\data_array.data0[6][62] ));
 sky130_fd_sc_hd__dfxtp_2 _12053_ (.CLK(clk),
    .D(_00861_),
    .Q(\data_array.data0[6][63] ));
 sky130_fd_sc_hd__dfxtp_2 _12054_ (.CLK(clk),
    .D(_00862_),
    .Q(\data_array.data1[14][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12055_ (.CLK(clk),
    .D(_00863_),
    .Q(\data_array.data1[14][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12056_ (.CLK(clk),
    .D(_00864_),
    .Q(\data_array.data1[14][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12057_ (.CLK(clk),
    .D(_00865_),
    .Q(\data_array.data1[14][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12058_ (.CLK(clk),
    .D(_00866_),
    .Q(\data_array.data1[14][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12059_ (.CLK(clk),
    .D(_00867_),
    .Q(\data_array.data1[14][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12060_ (.CLK(clk),
    .D(_00868_),
    .Q(\data_array.data1[14][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12061_ (.CLK(clk),
    .D(_00869_),
    .Q(\data_array.data1[14][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12062_ (.CLK(clk),
    .D(_00870_),
    .Q(\data_array.data1[14][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12063_ (.CLK(clk),
    .D(_00871_),
    .Q(\data_array.data1[14][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12064_ (.CLK(clk),
    .D(_00872_),
    .Q(\data_array.data1[14][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12065_ (.CLK(clk),
    .D(_00873_),
    .Q(\data_array.data1[14][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12066_ (.CLK(clk),
    .D(_00874_),
    .Q(\data_array.data1[14][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12067_ (.CLK(clk),
    .D(_00875_),
    .Q(\data_array.data1[14][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12068_ (.CLK(clk),
    .D(_00876_),
    .Q(\data_array.data1[14][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12069_ (.CLK(clk),
    .D(_00877_),
    .Q(\data_array.data1[14][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12070_ (.CLK(clk),
    .D(_00878_),
    .Q(\data_array.data1[14][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12071_ (.CLK(clk),
    .D(_00879_),
    .Q(\data_array.data1[14][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12072_ (.CLK(clk),
    .D(_00880_),
    .Q(\data_array.data1[14][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12073_ (.CLK(clk),
    .D(_00881_),
    .Q(\data_array.data1[14][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12074_ (.CLK(clk),
    .D(_00882_),
    .Q(\data_array.data1[14][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12075_ (.CLK(clk),
    .D(_00883_),
    .Q(\data_array.data1[14][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12076_ (.CLK(clk),
    .D(_00884_),
    .Q(\data_array.data1[14][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12077_ (.CLK(clk),
    .D(_00885_),
    .Q(\data_array.data1[14][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12078_ (.CLK(clk),
    .D(_00886_),
    .Q(\data_array.data1[14][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12079_ (.CLK(clk),
    .D(_00887_),
    .Q(\data_array.data1[14][25] ));
 sky130_fd_sc_hd__dfxtp_2 _12080_ (.CLK(clk),
    .D(_00888_),
    .Q(\data_array.data1[14][26] ));
 sky130_fd_sc_hd__dfxtp_2 _12081_ (.CLK(clk),
    .D(_00889_),
    .Q(\data_array.data1[14][27] ));
 sky130_fd_sc_hd__dfxtp_2 _12082_ (.CLK(clk),
    .D(_00890_),
    .Q(\data_array.data1[14][28] ));
 sky130_fd_sc_hd__dfxtp_2 _12083_ (.CLK(clk),
    .D(_00891_),
    .Q(\data_array.data1[14][29] ));
 sky130_fd_sc_hd__dfxtp_2 _12084_ (.CLK(clk),
    .D(_00892_),
    .Q(\data_array.data1[14][30] ));
 sky130_fd_sc_hd__dfxtp_2 _12085_ (.CLK(clk),
    .D(_00893_),
    .Q(\data_array.data1[14][31] ));
 sky130_fd_sc_hd__dfxtp_2 _12086_ (.CLK(clk),
    .D(_00894_),
    .Q(\data_array.data1[14][32] ));
 sky130_fd_sc_hd__dfxtp_2 _12087_ (.CLK(clk),
    .D(_00895_),
    .Q(\data_array.data1[14][33] ));
 sky130_fd_sc_hd__dfxtp_2 _12088_ (.CLK(clk),
    .D(_00896_),
    .Q(\data_array.data1[14][34] ));
 sky130_fd_sc_hd__dfxtp_2 _12089_ (.CLK(clk),
    .D(_00897_),
    .Q(\data_array.data1[14][35] ));
 sky130_fd_sc_hd__dfxtp_2 _12090_ (.CLK(clk),
    .D(_00898_),
    .Q(\data_array.data1[14][36] ));
 sky130_fd_sc_hd__dfxtp_2 _12091_ (.CLK(clk),
    .D(_00899_),
    .Q(\data_array.data1[14][37] ));
 sky130_fd_sc_hd__dfxtp_2 _12092_ (.CLK(clk),
    .D(_00900_),
    .Q(\data_array.data1[14][38] ));
 sky130_fd_sc_hd__dfxtp_2 _12093_ (.CLK(clk),
    .D(_00901_),
    .Q(\data_array.data1[14][39] ));
 sky130_fd_sc_hd__dfxtp_2 _12094_ (.CLK(clk),
    .D(_00902_),
    .Q(\data_array.data1[14][40] ));
 sky130_fd_sc_hd__dfxtp_2 _12095_ (.CLK(clk),
    .D(_00903_),
    .Q(\data_array.data1[14][41] ));
 sky130_fd_sc_hd__dfxtp_2 _12096_ (.CLK(clk),
    .D(_00904_),
    .Q(\data_array.data1[14][42] ));
 sky130_fd_sc_hd__dfxtp_2 _12097_ (.CLK(clk),
    .D(_00905_),
    .Q(\data_array.data1[14][43] ));
 sky130_fd_sc_hd__dfxtp_2 _12098_ (.CLK(clk),
    .D(_00906_),
    .Q(\data_array.data1[14][44] ));
 sky130_fd_sc_hd__dfxtp_2 _12099_ (.CLK(clk),
    .D(_00907_),
    .Q(\data_array.data1[14][45] ));
 sky130_fd_sc_hd__dfxtp_2 _12100_ (.CLK(clk),
    .D(_00908_),
    .Q(\data_array.data1[14][46] ));
 sky130_fd_sc_hd__dfxtp_2 _12101_ (.CLK(clk),
    .D(_00909_),
    .Q(\data_array.data1[14][47] ));
 sky130_fd_sc_hd__dfxtp_2 _12102_ (.CLK(clk),
    .D(_00910_),
    .Q(\data_array.data1[14][48] ));
 sky130_fd_sc_hd__dfxtp_2 _12103_ (.CLK(clk),
    .D(_00911_),
    .Q(\data_array.data1[14][49] ));
 sky130_fd_sc_hd__dfxtp_2 _12104_ (.CLK(clk),
    .D(_00912_),
    .Q(\data_array.data1[14][50] ));
 sky130_fd_sc_hd__dfxtp_2 _12105_ (.CLK(clk),
    .D(_00913_),
    .Q(\data_array.data1[14][51] ));
 sky130_fd_sc_hd__dfxtp_2 _12106_ (.CLK(clk),
    .D(_00914_),
    .Q(\data_array.data1[14][52] ));
 sky130_fd_sc_hd__dfxtp_2 _12107_ (.CLK(clk),
    .D(_00915_),
    .Q(\data_array.data1[14][53] ));
 sky130_fd_sc_hd__dfxtp_2 _12108_ (.CLK(clk),
    .D(_00916_),
    .Q(\data_array.data1[14][54] ));
 sky130_fd_sc_hd__dfxtp_2 _12109_ (.CLK(clk),
    .D(_00917_),
    .Q(\data_array.data1[14][55] ));
 sky130_fd_sc_hd__dfxtp_2 _12110_ (.CLK(clk),
    .D(_00918_),
    .Q(\data_array.data1[14][56] ));
 sky130_fd_sc_hd__dfxtp_2 _12111_ (.CLK(clk),
    .D(_00919_),
    .Q(\data_array.data1[14][57] ));
 sky130_fd_sc_hd__dfxtp_2 _12112_ (.CLK(clk),
    .D(_00920_),
    .Q(\data_array.data1[14][58] ));
 sky130_fd_sc_hd__dfxtp_2 _12113_ (.CLK(clk),
    .D(_00921_),
    .Q(\data_array.data1[14][59] ));
 sky130_fd_sc_hd__dfxtp_2 _12114_ (.CLK(clk),
    .D(_00922_),
    .Q(\data_array.data1[14][60] ));
 sky130_fd_sc_hd__dfxtp_2 _12115_ (.CLK(clk),
    .D(_00923_),
    .Q(\data_array.data1[14][61] ));
 sky130_fd_sc_hd__dfxtp_2 _12116_ (.CLK(clk),
    .D(_00924_),
    .Q(\data_array.data1[14][62] ));
 sky130_fd_sc_hd__dfxtp_2 _12117_ (.CLK(clk),
    .D(_00925_),
    .Q(\data_array.data1[14][63] ));
 sky130_fd_sc_hd__dfxtp_2 _12118_ (.CLK(clk),
    .D(_00926_),
    .Q(\tag_array.tag0[12][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12119_ (.CLK(clk),
    .D(_00927_),
    .Q(\tag_array.tag0[12][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12120_ (.CLK(clk),
    .D(_00928_),
    .Q(\tag_array.tag0[12][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12121_ (.CLK(clk),
    .D(_00929_),
    .Q(\tag_array.tag0[12][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12122_ (.CLK(clk),
    .D(_00930_),
    .Q(\tag_array.tag0[12][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12123_ (.CLK(clk),
    .D(_00931_),
    .Q(\tag_array.tag0[12][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12124_ (.CLK(clk),
    .D(_00932_),
    .Q(\tag_array.tag0[12][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12125_ (.CLK(clk),
    .D(_00933_),
    .Q(\tag_array.tag0[12][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12126_ (.CLK(clk),
    .D(_00934_),
    .Q(\tag_array.tag0[12][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12127_ (.CLK(clk),
    .D(_00935_),
    .Q(\tag_array.tag0[12][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12128_ (.CLK(clk),
    .D(_00936_),
    .Q(\tag_array.tag0[12][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12129_ (.CLK(clk),
    .D(_00937_),
    .Q(\tag_array.tag0[12][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12130_ (.CLK(clk),
    .D(_00938_),
    .Q(\tag_array.tag0[12][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12131_ (.CLK(clk),
    .D(_00939_),
    .Q(\tag_array.tag0[12][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12132_ (.CLK(clk),
    .D(_00940_),
    .Q(\tag_array.tag0[12][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12133_ (.CLK(clk),
    .D(_00941_),
    .Q(\tag_array.tag0[12][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12134_ (.CLK(clk),
    .D(_00942_),
    .Q(\tag_array.tag0[12][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12135_ (.CLK(clk),
    .D(_00943_),
    .Q(\tag_array.tag0[12][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12136_ (.CLK(clk),
    .D(_00944_),
    .Q(\tag_array.tag0[12][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12137_ (.CLK(clk),
    .D(_00945_),
    .Q(\tag_array.tag0[12][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12138_ (.CLK(clk),
    .D(_00946_),
    .Q(\tag_array.tag0[12][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12139_ (.CLK(clk),
    .D(_00947_),
    .Q(\tag_array.tag0[12][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12140_ (.CLK(clk),
    .D(_00948_),
    .Q(\tag_array.tag0[12][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12141_ (.CLK(clk),
    .D(_00949_),
    .Q(\tag_array.tag0[12][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12142_ (.CLK(clk),
    .D(_00950_),
    .Q(\tag_array.tag0[12][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12143_ (.CLK(clk),
    .D(_00951_),
    .Q(\tag_array.tag0[13][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12144_ (.CLK(clk),
    .D(_00952_),
    .Q(\tag_array.tag0[13][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12145_ (.CLK(clk),
    .D(_00953_),
    .Q(\tag_array.tag0[13][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12146_ (.CLK(clk),
    .D(_00954_),
    .Q(\tag_array.tag0[13][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12147_ (.CLK(clk),
    .D(_00955_),
    .Q(\tag_array.tag0[13][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12148_ (.CLK(clk),
    .D(_00956_),
    .Q(\tag_array.tag0[13][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12149_ (.CLK(clk),
    .D(_00957_),
    .Q(\tag_array.tag0[13][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12150_ (.CLK(clk),
    .D(_00958_),
    .Q(\tag_array.tag0[13][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12151_ (.CLK(clk),
    .D(_00959_),
    .Q(\tag_array.tag0[13][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12152_ (.CLK(clk),
    .D(_00960_),
    .Q(\tag_array.tag0[13][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12153_ (.CLK(clk),
    .D(_00961_),
    .Q(\tag_array.tag0[13][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12154_ (.CLK(clk),
    .D(_00962_),
    .Q(\tag_array.tag0[13][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12155_ (.CLK(clk),
    .D(_00963_),
    .Q(\tag_array.tag0[13][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12156_ (.CLK(clk),
    .D(_00964_),
    .Q(\tag_array.tag0[13][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12157_ (.CLK(clk),
    .D(_00965_),
    .Q(\tag_array.tag0[13][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12158_ (.CLK(clk),
    .D(_00966_),
    .Q(\tag_array.tag0[13][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12159_ (.CLK(clk),
    .D(_00967_),
    .Q(\tag_array.tag0[13][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12160_ (.CLK(clk),
    .D(_00968_),
    .Q(\tag_array.tag0[13][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12161_ (.CLK(clk),
    .D(_00969_),
    .Q(\tag_array.tag0[13][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12162_ (.CLK(clk),
    .D(_00970_),
    .Q(\tag_array.tag0[13][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12163_ (.CLK(clk),
    .D(_00971_),
    .Q(\tag_array.tag0[13][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12164_ (.CLK(clk),
    .D(_00972_),
    .Q(\tag_array.tag0[13][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12165_ (.CLK(clk),
    .D(_00973_),
    .Q(\tag_array.tag0[13][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12166_ (.CLK(clk),
    .D(_00974_),
    .Q(\tag_array.tag0[13][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12167_ (.CLK(clk),
    .D(_00975_),
    .Q(\tag_array.tag0[13][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12168_ (.CLK(clk),
    .D(_00976_),
    .Q(\tag_array.tag0[14][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12169_ (.CLK(clk),
    .D(_00977_),
    .Q(\tag_array.tag0[14][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12170_ (.CLK(clk),
    .D(_00978_),
    .Q(\tag_array.tag0[14][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12171_ (.CLK(clk),
    .D(_00979_),
    .Q(\tag_array.tag0[14][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12172_ (.CLK(clk),
    .D(_00980_),
    .Q(\tag_array.tag0[14][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12173_ (.CLK(clk),
    .D(_00981_),
    .Q(\tag_array.tag0[14][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12174_ (.CLK(clk),
    .D(_00982_),
    .Q(\tag_array.tag0[14][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12175_ (.CLK(clk),
    .D(_00983_),
    .Q(\tag_array.tag0[14][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12176_ (.CLK(clk),
    .D(_00984_),
    .Q(\tag_array.tag0[14][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12177_ (.CLK(clk),
    .D(_00985_),
    .Q(\tag_array.tag0[14][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12178_ (.CLK(clk),
    .D(_00986_),
    .Q(\tag_array.tag0[14][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12179_ (.CLK(clk),
    .D(_00987_),
    .Q(\tag_array.tag0[14][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12180_ (.CLK(clk),
    .D(_00988_),
    .Q(\tag_array.tag0[14][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12181_ (.CLK(clk),
    .D(_00989_),
    .Q(\tag_array.tag0[14][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12182_ (.CLK(clk),
    .D(_00990_),
    .Q(\tag_array.tag0[14][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12183_ (.CLK(clk),
    .D(_00991_),
    .Q(\tag_array.tag0[14][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12184_ (.CLK(clk),
    .D(_00992_),
    .Q(\tag_array.tag0[14][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12185_ (.CLK(clk),
    .D(_00993_),
    .Q(\tag_array.tag0[14][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12186_ (.CLK(clk),
    .D(_00994_),
    .Q(\tag_array.tag0[14][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12187_ (.CLK(clk),
    .D(_00995_),
    .Q(\tag_array.tag0[14][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12188_ (.CLK(clk),
    .D(_00996_),
    .Q(\tag_array.tag0[14][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12189_ (.CLK(clk),
    .D(_00997_),
    .Q(\tag_array.tag0[14][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12190_ (.CLK(clk),
    .D(_00998_),
    .Q(\tag_array.tag0[14][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12191_ (.CLK(clk),
    .D(_00999_),
    .Q(\tag_array.tag0[14][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12192_ (.CLK(clk),
    .D(_01000_),
    .Q(\tag_array.tag0[14][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12193_ (.CLK(clk),
    .D(_00131_),
    .Q(\fsm.tag_out0[0] ));
 sky130_fd_sc_hd__dfxtp_2 _12194_ (.CLK(clk),
    .D(_00142_),
    .Q(\fsm.tag_out0[1] ));
 sky130_fd_sc_hd__dfxtp_2 _12195_ (.CLK(clk),
    .D(_00148_),
    .Q(\fsm.tag_out0[2] ));
 sky130_fd_sc_hd__dfxtp_2 _12196_ (.CLK(clk),
    .D(_00149_),
    .Q(\fsm.tag_out0[3] ));
 sky130_fd_sc_hd__dfxtp_2 _12197_ (.CLK(clk),
    .D(_00150_),
    .Q(\fsm.tag_out0[4] ));
 sky130_fd_sc_hd__dfxtp_2 _12198_ (.CLK(clk),
    .D(_00151_),
    .Q(\fsm.tag_out0[5] ));
 sky130_fd_sc_hd__dfxtp_2 _12199_ (.CLK(clk),
    .D(_00152_),
    .Q(\fsm.tag_out0[6] ));
 sky130_fd_sc_hd__dfxtp_2 _12200_ (.CLK(clk),
    .D(_00153_),
    .Q(\fsm.tag_out0[7] ));
 sky130_fd_sc_hd__dfxtp_2 _12201_ (.CLK(clk),
    .D(_00154_),
    .Q(\fsm.tag_out0[8] ));
 sky130_fd_sc_hd__dfxtp_2 _12202_ (.CLK(clk),
    .D(_00155_),
    .Q(\fsm.tag_out0[9] ));
 sky130_fd_sc_hd__dfxtp_2 _12203_ (.CLK(clk),
    .D(_00132_),
    .Q(\fsm.tag_out0[10] ));
 sky130_fd_sc_hd__dfxtp_2 _12204_ (.CLK(clk),
    .D(_00133_),
    .Q(\fsm.tag_out0[11] ));
 sky130_fd_sc_hd__dfxtp_2 _12205_ (.CLK(clk),
    .D(_00134_),
    .Q(\fsm.tag_out0[12] ));
 sky130_fd_sc_hd__dfxtp_2 _12206_ (.CLK(clk),
    .D(_00135_),
    .Q(\fsm.tag_out0[13] ));
 sky130_fd_sc_hd__dfxtp_2 _12207_ (.CLK(clk),
    .D(_00136_),
    .Q(\fsm.tag_out0[14] ));
 sky130_fd_sc_hd__dfxtp_2 _12208_ (.CLK(clk),
    .D(_00137_),
    .Q(\fsm.tag_out0[15] ));
 sky130_fd_sc_hd__dfxtp_2 _12209_ (.CLK(clk),
    .D(_00138_),
    .Q(\fsm.tag_out0[16] ));
 sky130_fd_sc_hd__dfxtp_2 _12210_ (.CLK(clk),
    .D(_00139_),
    .Q(\fsm.tag_out0[17] ));
 sky130_fd_sc_hd__dfxtp_2 _12211_ (.CLK(clk),
    .D(_00140_),
    .Q(\fsm.tag_out0[18] ));
 sky130_fd_sc_hd__dfxtp_2 _12212_ (.CLK(clk),
    .D(_00141_),
    .Q(\fsm.tag_out0[19] ));
 sky130_fd_sc_hd__dfxtp_2 _12213_ (.CLK(clk),
    .D(_00143_),
    .Q(\fsm.tag_out0[20] ));
 sky130_fd_sc_hd__dfxtp_2 _12214_ (.CLK(clk),
    .D(_00144_),
    .Q(\fsm.tag_out0[21] ));
 sky130_fd_sc_hd__dfxtp_2 _12215_ (.CLK(clk),
    .D(_00145_),
    .Q(\fsm.tag_out0[22] ));
 sky130_fd_sc_hd__dfxtp_2 _12216_ (.CLK(clk),
    .D(_00146_),
    .Q(\fsm.tag_out0[23] ));
 sky130_fd_sc_hd__dfxtp_2 _12217_ (.CLK(clk),
    .D(_00147_),
    .Q(\fsm.tag_out0[24] ));
 sky130_fd_sc_hd__dfxtp_2 _12218_ (.CLK(clk),
    .D(_00156_),
    .Q(\fsm.tag_out1[0] ));
 sky130_fd_sc_hd__dfxtp_2 _12219_ (.CLK(clk),
    .D(_00167_),
    .Q(\fsm.tag_out1[1] ));
 sky130_fd_sc_hd__dfxtp_2 _12220_ (.CLK(clk),
    .D(_00173_),
    .Q(\fsm.tag_out1[2] ));
 sky130_fd_sc_hd__dfxtp_2 _12221_ (.CLK(clk),
    .D(_00174_),
    .Q(\fsm.tag_out1[3] ));
 sky130_fd_sc_hd__dfxtp_2 _12222_ (.CLK(clk),
    .D(_00175_),
    .Q(\fsm.tag_out1[4] ));
 sky130_fd_sc_hd__dfxtp_2 _12223_ (.CLK(clk),
    .D(_00176_),
    .Q(\fsm.tag_out1[5] ));
 sky130_fd_sc_hd__dfxtp_2 _12224_ (.CLK(clk),
    .D(_00177_),
    .Q(\fsm.tag_out1[6] ));
 sky130_fd_sc_hd__dfxtp_2 _12225_ (.CLK(clk),
    .D(_00178_),
    .Q(\fsm.tag_out1[7] ));
 sky130_fd_sc_hd__dfxtp_2 _12226_ (.CLK(clk),
    .D(_00179_),
    .Q(\fsm.tag_out1[8] ));
 sky130_fd_sc_hd__dfxtp_2 _12227_ (.CLK(clk),
    .D(_00180_),
    .Q(\fsm.tag_out1[9] ));
 sky130_fd_sc_hd__dfxtp_2 _12228_ (.CLK(clk),
    .D(_00157_),
    .Q(\fsm.tag_out1[10] ));
 sky130_fd_sc_hd__dfxtp_2 _12229_ (.CLK(clk),
    .D(_00158_),
    .Q(\fsm.tag_out1[11] ));
 sky130_fd_sc_hd__dfxtp_2 _12230_ (.CLK(clk),
    .D(_00159_),
    .Q(\fsm.tag_out1[12] ));
 sky130_fd_sc_hd__dfxtp_2 _12231_ (.CLK(clk),
    .D(_00160_),
    .Q(\fsm.tag_out1[13] ));
 sky130_fd_sc_hd__dfxtp_2 _12232_ (.CLK(clk),
    .D(_00161_),
    .Q(\fsm.tag_out1[14] ));
 sky130_fd_sc_hd__dfxtp_2 _12233_ (.CLK(clk),
    .D(_00162_),
    .Q(\fsm.tag_out1[15] ));
 sky130_fd_sc_hd__dfxtp_2 _12234_ (.CLK(clk),
    .D(_00163_),
    .Q(\fsm.tag_out1[16] ));
 sky130_fd_sc_hd__dfxtp_2 _12235_ (.CLK(clk),
    .D(_00164_),
    .Q(\fsm.tag_out1[17] ));
 sky130_fd_sc_hd__dfxtp_2 _12236_ (.CLK(clk),
    .D(_00165_),
    .Q(\fsm.tag_out1[18] ));
 sky130_fd_sc_hd__dfxtp_2 _12237_ (.CLK(clk),
    .D(_00166_),
    .Q(\fsm.tag_out1[19] ));
 sky130_fd_sc_hd__dfxtp_2 _12238_ (.CLK(clk),
    .D(_00168_),
    .Q(\fsm.tag_out1[20] ));
 sky130_fd_sc_hd__dfxtp_2 _12239_ (.CLK(clk),
    .D(_00169_),
    .Q(\fsm.tag_out1[21] ));
 sky130_fd_sc_hd__dfxtp_2 _12240_ (.CLK(clk),
    .D(_00170_),
    .Q(\fsm.tag_out1[22] ));
 sky130_fd_sc_hd__dfxtp_2 _12241_ (.CLK(clk),
    .D(_00171_),
    .Q(\fsm.tag_out1[23] ));
 sky130_fd_sc_hd__dfxtp_2 _12242_ (.CLK(clk),
    .D(_00172_),
    .Q(\fsm.tag_out1[24] ));
 sky130_fd_sc_hd__dfxtp_2 _12243_ (.CLK(clk),
    .D(_01001_),
    .Q(\tag_array.tag1[14][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12244_ (.CLK(clk),
    .D(_01002_),
    .Q(\tag_array.tag1[14][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12245_ (.CLK(clk),
    .D(_01003_),
    .Q(\tag_array.tag1[14][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12246_ (.CLK(clk),
    .D(_01004_),
    .Q(\tag_array.tag1[14][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12247_ (.CLK(clk),
    .D(_01005_),
    .Q(\tag_array.tag1[14][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12248_ (.CLK(clk),
    .D(_01006_),
    .Q(\tag_array.tag1[14][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12249_ (.CLK(clk),
    .D(_01007_),
    .Q(\tag_array.tag1[14][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12250_ (.CLK(clk),
    .D(_01008_),
    .Q(\tag_array.tag1[14][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12251_ (.CLK(clk),
    .D(_01009_),
    .Q(\tag_array.tag1[14][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12252_ (.CLK(clk),
    .D(_01010_),
    .Q(\tag_array.tag1[14][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12253_ (.CLK(clk),
    .D(_01011_),
    .Q(\tag_array.tag1[14][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12254_ (.CLK(clk),
    .D(_01012_),
    .Q(\tag_array.tag1[14][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12255_ (.CLK(clk),
    .D(_01013_),
    .Q(\tag_array.tag1[14][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12256_ (.CLK(clk),
    .D(_01014_),
    .Q(\tag_array.tag1[14][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12257_ (.CLK(clk),
    .D(_01015_),
    .Q(\tag_array.tag1[14][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12258_ (.CLK(clk),
    .D(_01016_),
    .Q(\tag_array.tag1[14][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12259_ (.CLK(clk),
    .D(_01017_),
    .Q(\tag_array.tag1[14][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12260_ (.CLK(clk),
    .D(_01018_),
    .Q(\tag_array.tag1[14][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12261_ (.CLK(clk),
    .D(_01019_),
    .Q(\tag_array.tag1[14][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12262_ (.CLK(clk),
    .D(_01020_),
    .Q(\tag_array.tag1[14][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12263_ (.CLK(clk),
    .D(_01021_),
    .Q(\tag_array.tag1[14][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12264_ (.CLK(clk),
    .D(_01022_),
    .Q(\tag_array.tag1[14][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12265_ (.CLK(clk),
    .D(_01023_),
    .Q(\tag_array.tag1[14][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12266_ (.CLK(clk),
    .D(_01024_),
    .Q(\tag_array.tag1[14][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12267_ (.CLK(clk),
    .D(_01025_),
    .Q(\tag_array.tag1[14][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12268_ (.CLK(clk),
    .D(_01026_),
    .Q(\tag_array.tag1[13][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12269_ (.CLK(clk),
    .D(_01027_),
    .Q(\tag_array.tag1[13][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12270_ (.CLK(clk),
    .D(_01028_),
    .Q(\tag_array.tag1[13][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12271_ (.CLK(clk),
    .D(_01029_),
    .Q(\tag_array.tag1[13][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12272_ (.CLK(clk),
    .D(_01030_),
    .Q(\tag_array.tag1[13][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12273_ (.CLK(clk),
    .D(_01031_),
    .Q(\tag_array.tag1[13][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12274_ (.CLK(clk),
    .D(_01032_),
    .Q(\tag_array.tag1[13][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12275_ (.CLK(clk),
    .D(_01033_),
    .Q(\tag_array.tag1[13][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12276_ (.CLK(clk),
    .D(_01034_),
    .Q(\tag_array.tag1[13][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12277_ (.CLK(clk),
    .D(_01035_),
    .Q(\tag_array.tag1[13][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12278_ (.CLK(clk),
    .D(_01036_),
    .Q(\tag_array.tag1[13][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12279_ (.CLK(clk),
    .D(_01037_),
    .Q(\tag_array.tag1[13][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12280_ (.CLK(clk),
    .D(_01038_),
    .Q(\tag_array.tag1[13][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12281_ (.CLK(clk),
    .D(_01039_),
    .Q(\tag_array.tag1[13][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12282_ (.CLK(clk),
    .D(_01040_),
    .Q(\tag_array.tag1[13][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12283_ (.CLK(clk),
    .D(_01041_),
    .Q(\tag_array.tag1[13][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12284_ (.CLK(clk),
    .D(_01042_),
    .Q(\tag_array.tag1[13][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12285_ (.CLK(clk),
    .D(_01043_),
    .Q(\tag_array.tag1[13][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12286_ (.CLK(clk),
    .D(_01044_),
    .Q(\tag_array.tag1[13][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12287_ (.CLK(clk),
    .D(_01045_),
    .Q(\tag_array.tag1[13][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12288_ (.CLK(clk),
    .D(_01046_),
    .Q(\tag_array.tag1[13][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12289_ (.CLK(clk),
    .D(_01047_),
    .Q(\tag_array.tag1[13][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12290_ (.CLK(clk),
    .D(_01048_),
    .Q(\tag_array.tag1[13][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12291_ (.CLK(clk),
    .D(_01049_),
    .Q(\tag_array.tag1[13][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12292_ (.CLK(clk),
    .D(_01050_),
    .Q(\tag_array.tag1[13][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12293_ (.CLK(clk),
    .D(_01051_),
    .Q(\tag_array.tag1[12][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12294_ (.CLK(clk),
    .D(_01052_),
    .Q(\tag_array.tag1[12][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12295_ (.CLK(clk),
    .D(_01053_),
    .Q(\tag_array.tag1[12][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12296_ (.CLK(clk),
    .D(_01054_),
    .Q(\tag_array.tag1[12][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12297_ (.CLK(clk),
    .D(_01055_),
    .Q(\tag_array.tag1[12][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12298_ (.CLK(clk),
    .D(_01056_),
    .Q(\tag_array.tag1[12][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12299_ (.CLK(clk),
    .D(_01057_),
    .Q(\tag_array.tag1[12][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12300_ (.CLK(clk),
    .D(_01058_),
    .Q(\tag_array.tag1[12][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12301_ (.CLK(clk),
    .D(_01059_),
    .Q(\tag_array.tag1[12][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12302_ (.CLK(clk),
    .D(_01060_),
    .Q(\tag_array.tag1[12][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12303_ (.CLK(clk),
    .D(_01061_),
    .Q(\tag_array.tag1[12][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12304_ (.CLK(clk),
    .D(_01062_),
    .Q(\tag_array.tag1[12][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12305_ (.CLK(clk),
    .D(_01063_),
    .Q(\tag_array.tag1[12][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12306_ (.CLK(clk),
    .D(_01064_),
    .Q(\tag_array.tag1[12][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12307_ (.CLK(clk),
    .D(_01065_),
    .Q(\tag_array.tag1[12][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12308_ (.CLK(clk),
    .D(_01066_),
    .Q(\tag_array.tag1[12][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12309_ (.CLK(clk),
    .D(_01067_),
    .Q(\tag_array.tag1[12][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12310_ (.CLK(clk),
    .D(_01068_),
    .Q(\tag_array.tag1[12][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12311_ (.CLK(clk),
    .D(_01069_),
    .Q(\tag_array.tag1[12][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12312_ (.CLK(clk),
    .D(_01070_),
    .Q(\tag_array.tag1[12][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12313_ (.CLK(clk),
    .D(_01071_),
    .Q(\tag_array.tag1[12][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12314_ (.CLK(clk),
    .D(_01072_),
    .Q(\tag_array.tag1[12][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12315_ (.CLK(clk),
    .D(_01073_),
    .Q(\tag_array.tag1[12][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12316_ (.CLK(clk),
    .D(_01074_),
    .Q(\tag_array.tag1[12][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12317_ (.CLK(clk),
    .D(_01075_),
    .Q(\tag_array.tag1[12][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12318_ (.CLK(clk),
    .D(_00000_),
    .Q(\data_array.rdata0[0] ));
 sky130_fd_sc_hd__dfxtp_2 _12319_ (.CLK(clk),
    .D(_00011_),
    .Q(\data_array.rdata0[1] ));
 sky130_fd_sc_hd__dfxtp_2 _12320_ (.CLK(clk),
    .D(_00022_),
    .Q(\data_array.rdata0[2] ));
 sky130_fd_sc_hd__dfxtp_2 _12321_ (.CLK(clk),
    .D(_00033_),
    .Q(\data_array.rdata0[3] ));
 sky130_fd_sc_hd__dfxtp_2 _12322_ (.CLK(clk),
    .D(_00044_),
    .Q(\data_array.rdata0[4] ));
 sky130_fd_sc_hd__dfxtp_2 _12323_ (.CLK(clk),
    .D(_00055_),
    .Q(\data_array.rdata0[5] ));
 sky130_fd_sc_hd__dfxtp_2 _12324_ (.CLK(clk),
    .D(_00060_),
    .Q(\data_array.rdata0[6] ));
 sky130_fd_sc_hd__dfxtp_2 _12325_ (.CLK(clk),
    .D(_00061_),
    .Q(\data_array.rdata0[7] ));
 sky130_fd_sc_hd__dfxtp_2 _12326_ (.CLK(clk),
    .D(_00062_),
    .Q(\data_array.rdata0[8] ));
 sky130_fd_sc_hd__dfxtp_2 _12327_ (.CLK(clk),
    .D(_00063_),
    .Q(\data_array.rdata0[9] ));
 sky130_fd_sc_hd__dfxtp_2 _12328_ (.CLK(clk),
    .D(_00001_),
    .Q(\data_array.rdata0[10] ));
 sky130_fd_sc_hd__dfxtp_2 _12329_ (.CLK(clk),
    .D(_00002_),
    .Q(\data_array.rdata0[11] ));
 sky130_fd_sc_hd__dfxtp_2 _12330_ (.CLK(clk),
    .D(_00003_),
    .Q(\data_array.rdata0[12] ));
 sky130_fd_sc_hd__dfxtp_2 _12331_ (.CLK(clk),
    .D(_00004_),
    .Q(\data_array.rdata0[13] ));
 sky130_fd_sc_hd__dfxtp_2 _12332_ (.CLK(clk),
    .D(_00005_),
    .Q(\data_array.rdata0[14] ));
 sky130_fd_sc_hd__dfxtp_2 _12333_ (.CLK(clk),
    .D(_00006_),
    .Q(\data_array.rdata0[15] ));
 sky130_fd_sc_hd__dfxtp_2 _12334_ (.CLK(clk),
    .D(_00007_),
    .Q(\data_array.rdata0[16] ));
 sky130_fd_sc_hd__dfxtp_2 _12335_ (.CLK(clk),
    .D(_00008_),
    .Q(\data_array.rdata0[17] ));
 sky130_fd_sc_hd__dfxtp_2 _12336_ (.CLK(clk),
    .D(_00009_),
    .Q(\data_array.rdata0[18] ));
 sky130_fd_sc_hd__dfxtp_2 _12337_ (.CLK(clk),
    .D(_00010_),
    .Q(\data_array.rdata0[19] ));
 sky130_fd_sc_hd__dfxtp_2 _12338_ (.CLK(clk),
    .D(_00012_),
    .Q(\data_array.rdata0[20] ));
 sky130_fd_sc_hd__dfxtp_2 _12339_ (.CLK(clk),
    .D(_00013_),
    .Q(\data_array.rdata0[21] ));
 sky130_fd_sc_hd__dfxtp_2 _12340_ (.CLK(clk),
    .D(_00014_),
    .Q(\data_array.rdata0[22] ));
 sky130_fd_sc_hd__dfxtp_2 _12341_ (.CLK(clk),
    .D(_00015_),
    .Q(\data_array.rdata0[23] ));
 sky130_fd_sc_hd__dfxtp_2 _12342_ (.CLK(clk),
    .D(_00016_),
    .Q(\data_array.rdata0[24] ));
 sky130_fd_sc_hd__dfxtp_2 _12343_ (.CLK(clk),
    .D(_00017_),
    .Q(\data_array.rdata0[25] ));
 sky130_fd_sc_hd__dfxtp_2 _12344_ (.CLK(clk),
    .D(_00018_),
    .Q(\data_array.rdata0[26] ));
 sky130_fd_sc_hd__dfxtp_2 _12345_ (.CLK(clk),
    .D(_00019_),
    .Q(\data_array.rdata0[27] ));
 sky130_fd_sc_hd__dfxtp_2 _12346_ (.CLK(clk),
    .D(_00020_),
    .Q(\data_array.rdata0[28] ));
 sky130_fd_sc_hd__dfxtp_2 _12347_ (.CLK(clk),
    .D(_00021_),
    .Q(\data_array.rdata0[29] ));
 sky130_fd_sc_hd__dfxtp_2 _12348_ (.CLK(clk),
    .D(_00023_),
    .Q(\data_array.rdata0[30] ));
 sky130_fd_sc_hd__dfxtp_2 _12349_ (.CLK(clk),
    .D(_00024_),
    .Q(\data_array.rdata0[31] ));
 sky130_fd_sc_hd__dfxtp_2 _12350_ (.CLK(clk),
    .D(_00025_),
    .Q(\data_array.rdata0[32] ));
 sky130_fd_sc_hd__dfxtp_2 _12351_ (.CLK(clk),
    .D(_00026_),
    .Q(\data_array.rdata0[33] ));
 sky130_fd_sc_hd__dfxtp_2 _12352_ (.CLK(clk),
    .D(_00027_),
    .Q(\data_array.rdata0[34] ));
 sky130_fd_sc_hd__dfxtp_2 _12353_ (.CLK(clk),
    .D(_00028_),
    .Q(\data_array.rdata0[35] ));
 sky130_fd_sc_hd__dfxtp_2 _12354_ (.CLK(clk),
    .D(_00029_),
    .Q(\data_array.rdata0[36] ));
 sky130_fd_sc_hd__dfxtp_2 _12355_ (.CLK(clk),
    .D(_00030_),
    .Q(\data_array.rdata0[37] ));
 sky130_fd_sc_hd__dfxtp_2 _12356_ (.CLK(clk),
    .D(_00031_),
    .Q(\data_array.rdata0[38] ));
 sky130_fd_sc_hd__dfxtp_2 _12357_ (.CLK(clk),
    .D(_00032_),
    .Q(\data_array.rdata0[39] ));
 sky130_fd_sc_hd__dfxtp_2 _12358_ (.CLK(clk),
    .D(_00034_),
    .Q(\data_array.rdata0[40] ));
 sky130_fd_sc_hd__dfxtp_2 _12359_ (.CLK(clk),
    .D(_00035_),
    .Q(\data_array.rdata0[41] ));
 sky130_fd_sc_hd__dfxtp_2 _12360_ (.CLK(clk),
    .D(_00036_),
    .Q(\data_array.rdata0[42] ));
 sky130_fd_sc_hd__dfxtp_2 _12361_ (.CLK(clk),
    .D(_00037_),
    .Q(\data_array.rdata0[43] ));
 sky130_fd_sc_hd__dfxtp_2 _12362_ (.CLK(clk),
    .D(_00038_),
    .Q(\data_array.rdata0[44] ));
 sky130_fd_sc_hd__dfxtp_2 _12363_ (.CLK(clk),
    .D(_00039_),
    .Q(\data_array.rdata0[45] ));
 sky130_fd_sc_hd__dfxtp_2 _12364_ (.CLK(clk),
    .D(_00040_),
    .Q(\data_array.rdata0[46] ));
 sky130_fd_sc_hd__dfxtp_2 _12365_ (.CLK(clk),
    .D(_00041_),
    .Q(\data_array.rdata0[47] ));
 sky130_fd_sc_hd__dfxtp_2 _12366_ (.CLK(clk),
    .D(_00042_),
    .Q(\data_array.rdata0[48] ));
 sky130_fd_sc_hd__dfxtp_2 _12367_ (.CLK(clk),
    .D(_00043_),
    .Q(\data_array.rdata0[49] ));
 sky130_fd_sc_hd__dfxtp_2 _12368_ (.CLK(clk),
    .D(_00045_),
    .Q(\data_array.rdata0[50] ));
 sky130_fd_sc_hd__dfxtp_2 _12369_ (.CLK(clk),
    .D(_00046_),
    .Q(\data_array.rdata0[51] ));
 sky130_fd_sc_hd__dfxtp_2 _12370_ (.CLK(clk),
    .D(_00047_),
    .Q(\data_array.rdata0[52] ));
 sky130_fd_sc_hd__dfxtp_2 _12371_ (.CLK(clk),
    .D(_00048_),
    .Q(\data_array.rdata0[53] ));
 sky130_fd_sc_hd__dfxtp_2 _12372_ (.CLK(clk),
    .D(_00049_),
    .Q(\data_array.rdata0[54] ));
 sky130_fd_sc_hd__dfxtp_2 _12373_ (.CLK(clk),
    .D(_00050_),
    .Q(\data_array.rdata0[55] ));
 sky130_fd_sc_hd__dfxtp_2 _12374_ (.CLK(clk),
    .D(_00051_),
    .Q(\data_array.rdata0[56] ));
 sky130_fd_sc_hd__dfxtp_2 _12375_ (.CLK(clk),
    .D(_00052_),
    .Q(\data_array.rdata0[57] ));
 sky130_fd_sc_hd__dfxtp_2 _12376_ (.CLK(clk),
    .D(_00053_),
    .Q(\data_array.rdata0[58] ));
 sky130_fd_sc_hd__dfxtp_2 _12377_ (.CLK(clk),
    .D(_00054_),
    .Q(\data_array.rdata0[59] ));
 sky130_fd_sc_hd__dfxtp_2 _12378_ (.CLK(clk),
    .D(_00056_),
    .Q(\data_array.rdata0[60] ));
 sky130_fd_sc_hd__dfxtp_2 _12379_ (.CLK(clk),
    .D(_00057_),
    .Q(\data_array.rdata0[61] ));
 sky130_fd_sc_hd__dfxtp_2 _12380_ (.CLK(clk),
    .D(_00058_),
    .Q(\data_array.rdata0[62] ));
 sky130_fd_sc_hd__dfxtp_2 _12381_ (.CLK(clk),
    .D(_00059_),
    .Q(\data_array.rdata0[63] ));
 sky130_fd_sc_hd__dfxtp_2 _12382_ (.CLK(clk),
    .D(_01076_),
    .Q(\data_array.data0[14][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12383_ (.CLK(clk),
    .D(_01077_),
    .Q(\data_array.data0[14][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12384_ (.CLK(clk),
    .D(_01078_),
    .Q(\data_array.data0[14][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12385_ (.CLK(clk),
    .D(_01079_),
    .Q(\data_array.data0[14][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12386_ (.CLK(clk),
    .D(_01080_),
    .Q(\data_array.data0[14][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12387_ (.CLK(clk),
    .D(_01081_),
    .Q(\data_array.data0[14][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12388_ (.CLK(clk),
    .D(_01082_),
    .Q(\data_array.data0[14][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12389_ (.CLK(clk),
    .D(_01083_),
    .Q(\data_array.data0[14][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12390_ (.CLK(clk),
    .D(_01084_),
    .Q(\data_array.data0[14][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12391_ (.CLK(clk),
    .D(_01085_),
    .Q(\data_array.data0[14][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12392_ (.CLK(clk),
    .D(_01086_),
    .Q(\data_array.data0[14][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12393_ (.CLK(clk),
    .D(_01087_),
    .Q(\data_array.data0[14][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12394_ (.CLK(clk),
    .D(_01088_),
    .Q(\data_array.data0[14][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12395_ (.CLK(clk),
    .D(_01089_),
    .Q(\data_array.data0[14][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12396_ (.CLK(clk),
    .D(_01090_),
    .Q(\data_array.data0[14][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12397_ (.CLK(clk),
    .D(_01091_),
    .Q(\data_array.data0[14][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12398_ (.CLK(clk),
    .D(_01092_),
    .Q(\data_array.data0[14][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12399_ (.CLK(clk),
    .D(_01093_),
    .Q(\data_array.data0[14][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12400_ (.CLK(clk),
    .D(_01094_),
    .Q(\data_array.data0[14][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12401_ (.CLK(clk),
    .D(_01095_),
    .Q(\data_array.data0[14][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12402_ (.CLK(clk),
    .D(_01096_),
    .Q(\data_array.data0[14][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12403_ (.CLK(clk),
    .D(_01097_),
    .Q(\data_array.data0[14][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12404_ (.CLK(clk),
    .D(_01098_),
    .Q(\data_array.data0[14][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12405_ (.CLK(clk),
    .D(_01099_),
    .Q(\data_array.data0[14][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12406_ (.CLK(clk),
    .D(_01100_),
    .Q(\data_array.data0[14][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12407_ (.CLK(clk),
    .D(_01101_),
    .Q(\data_array.data0[14][25] ));
 sky130_fd_sc_hd__dfxtp_2 _12408_ (.CLK(clk),
    .D(_01102_),
    .Q(\data_array.data0[14][26] ));
 sky130_fd_sc_hd__dfxtp_2 _12409_ (.CLK(clk),
    .D(_01103_),
    .Q(\data_array.data0[14][27] ));
 sky130_fd_sc_hd__dfxtp_2 _12410_ (.CLK(clk),
    .D(_01104_),
    .Q(\data_array.data0[14][28] ));
 sky130_fd_sc_hd__dfxtp_2 _12411_ (.CLK(clk),
    .D(_01105_),
    .Q(\data_array.data0[14][29] ));
 sky130_fd_sc_hd__dfxtp_2 _12412_ (.CLK(clk),
    .D(_01106_),
    .Q(\data_array.data0[14][30] ));
 sky130_fd_sc_hd__dfxtp_2 _12413_ (.CLK(clk),
    .D(_01107_),
    .Q(\data_array.data0[14][31] ));
 sky130_fd_sc_hd__dfxtp_2 _12414_ (.CLK(clk),
    .D(_01108_),
    .Q(\data_array.data0[14][32] ));
 sky130_fd_sc_hd__dfxtp_2 _12415_ (.CLK(clk),
    .D(_01109_),
    .Q(\data_array.data0[14][33] ));
 sky130_fd_sc_hd__dfxtp_2 _12416_ (.CLK(clk),
    .D(_01110_),
    .Q(\data_array.data0[14][34] ));
 sky130_fd_sc_hd__dfxtp_2 _12417_ (.CLK(clk),
    .D(_01111_),
    .Q(\data_array.data0[14][35] ));
 sky130_fd_sc_hd__dfxtp_2 _12418_ (.CLK(clk),
    .D(_01112_),
    .Q(\data_array.data0[14][36] ));
 sky130_fd_sc_hd__dfxtp_2 _12419_ (.CLK(clk),
    .D(_01113_),
    .Q(\data_array.data0[14][37] ));
 sky130_fd_sc_hd__dfxtp_2 _12420_ (.CLK(clk),
    .D(_01114_),
    .Q(\data_array.data0[14][38] ));
 sky130_fd_sc_hd__dfxtp_2 _12421_ (.CLK(clk),
    .D(_01115_),
    .Q(\data_array.data0[14][39] ));
 sky130_fd_sc_hd__dfxtp_2 _12422_ (.CLK(clk),
    .D(_01116_),
    .Q(\data_array.data0[14][40] ));
 sky130_fd_sc_hd__dfxtp_2 _12423_ (.CLK(clk),
    .D(_01117_),
    .Q(\data_array.data0[14][41] ));
 sky130_fd_sc_hd__dfxtp_2 _12424_ (.CLK(clk),
    .D(_01118_),
    .Q(\data_array.data0[14][42] ));
 sky130_fd_sc_hd__dfxtp_2 _12425_ (.CLK(clk),
    .D(_01119_),
    .Q(\data_array.data0[14][43] ));
 sky130_fd_sc_hd__dfxtp_2 _12426_ (.CLK(clk),
    .D(_01120_),
    .Q(\data_array.data0[14][44] ));
 sky130_fd_sc_hd__dfxtp_2 _12427_ (.CLK(clk),
    .D(_01121_),
    .Q(\data_array.data0[14][45] ));
 sky130_fd_sc_hd__dfxtp_2 _12428_ (.CLK(clk),
    .D(_01122_),
    .Q(\data_array.data0[14][46] ));
 sky130_fd_sc_hd__dfxtp_2 _12429_ (.CLK(clk),
    .D(_01123_),
    .Q(\data_array.data0[14][47] ));
 sky130_fd_sc_hd__dfxtp_2 _12430_ (.CLK(clk),
    .D(_01124_),
    .Q(\data_array.data0[14][48] ));
 sky130_fd_sc_hd__dfxtp_2 _12431_ (.CLK(clk),
    .D(_01125_),
    .Q(\data_array.data0[14][49] ));
 sky130_fd_sc_hd__dfxtp_2 _12432_ (.CLK(clk),
    .D(_01126_),
    .Q(\data_array.data0[14][50] ));
 sky130_fd_sc_hd__dfxtp_2 _12433_ (.CLK(clk),
    .D(_01127_),
    .Q(\data_array.data0[14][51] ));
 sky130_fd_sc_hd__dfxtp_2 _12434_ (.CLK(clk),
    .D(_01128_),
    .Q(\data_array.data0[14][52] ));
 sky130_fd_sc_hd__dfxtp_2 _12435_ (.CLK(clk),
    .D(_01129_),
    .Q(\data_array.data0[14][53] ));
 sky130_fd_sc_hd__dfxtp_2 _12436_ (.CLK(clk),
    .D(_01130_),
    .Q(\data_array.data0[14][54] ));
 sky130_fd_sc_hd__dfxtp_2 _12437_ (.CLK(clk),
    .D(_01131_),
    .Q(\data_array.data0[14][55] ));
 sky130_fd_sc_hd__dfxtp_2 _12438_ (.CLK(clk),
    .D(_01132_),
    .Q(\data_array.data0[14][56] ));
 sky130_fd_sc_hd__dfxtp_2 _12439_ (.CLK(clk),
    .D(_01133_),
    .Q(\data_array.data0[14][57] ));
 sky130_fd_sc_hd__dfxtp_2 _12440_ (.CLK(clk),
    .D(_01134_),
    .Q(\data_array.data0[14][58] ));
 sky130_fd_sc_hd__dfxtp_2 _12441_ (.CLK(clk),
    .D(_01135_),
    .Q(\data_array.data0[14][59] ));
 sky130_fd_sc_hd__dfxtp_2 _12442_ (.CLK(clk),
    .D(_01136_),
    .Q(\data_array.data0[14][60] ));
 sky130_fd_sc_hd__dfxtp_2 _12443_ (.CLK(clk),
    .D(_01137_),
    .Q(\data_array.data0[14][61] ));
 sky130_fd_sc_hd__dfxtp_2 _12444_ (.CLK(clk),
    .D(_01138_),
    .Q(\data_array.data0[14][62] ));
 sky130_fd_sc_hd__dfxtp_2 _12445_ (.CLK(clk),
    .D(_01139_),
    .Q(\data_array.data0[14][63] ));
 sky130_fd_sc_hd__dfxtp_2 _12446_ (.CLK(clk),
    .D(_01140_),
    .Q(\lru_array.lru_mem[6] ));
 sky130_fd_sc_hd__dfxtp_2 _12447_ (.CLK(clk),
    .D(_01141_),
    .Q(\lru_array.lru_mem[7] ));
 sky130_fd_sc_hd__dfxtp_2 _12448_ (.CLK(clk),
    .D(_01142_),
    .Q(\data_array.data1[9][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12449_ (.CLK(clk),
    .D(_01143_),
    .Q(\data_array.data1[9][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12450_ (.CLK(clk),
    .D(_01144_),
    .Q(\data_array.data1[9][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12451_ (.CLK(clk),
    .D(_01145_),
    .Q(\data_array.data1[9][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12452_ (.CLK(clk),
    .D(_01146_),
    .Q(\data_array.data1[9][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12453_ (.CLK(clk),
    .D(_01147_),
    .Q(\data_array.data1[9][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12454_ (.CLK(clk),
    .D(_01148_),
    .Q(\data_array.data1[9][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12455_ (.CLK(clk),
    .D(_01149_),
    .Q(\data_array.data1[9][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12456_ (.CLK(clk),
    .D(_01150_),
    .Q(\data_array.data1[9][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12457_ (.CLK(clk),
    .D(_01151_),
    .Q(\data_array.data1[9][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12458_ (.CLK(clk),
    .D(_01152_),
    .Q(\data_array.data1[9][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12459_ (.CLK(clk),
    .D(_01153_),
    .Q(\data_array.data1[9][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12460_ (.CLK(clk),
    .D(_01154_),
    .Q(\data_array.data1[9][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12461_ (.CLK(clk),
    .D(_01155_),
    .Q(\data_array.data1[9][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12462_ (.CLK(clk),
    .D(_01156_),
    .Q(\data_array.data1[9][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12463_ (.CLK(clk),
    .D(_01157_),
    .Q(\data_array.data1[9][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12464_ (.CLK(clk),
    .D(_01158_),
    .Q(\data_array.data1[9][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12465_ (.CLK(clk),
    .D(_01159_),
    .Q(\data_array.data1[9][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12466_ (.CLK(clk),
    .D(_01160_),
    .Q(\data_array.data1[9][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12467_ (.CLK(clk),
    .D(_01161_),
    .Q(\data_array.data1[9][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12468_ (.CLK(clk),
    .D(_01162_),
    .Q(\data_array.data1[9][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12469_ (.CLK(clk),
    .D(_01163_),
    .Q(\data_array.data1[9][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12470_ (.CLK(clk),
    .D(_01164_),
    .Q(\data_array.data1[9][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12471_ (.CLK(clk),
    .D(_01165_),
    .Q(\data_array.data1[9][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12472_ (.CLK(clk),
    .D(_01166_),
    .Q(\data_array.data1[9][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12473_ (.CLK(clk),
    .D(_01167_),
    .Q(\data_array.data1[9][25] ));
 sky130_fd_sc_hd__dfxtp_2 _12474_ (.CLK(clk),
    .D(_01168_),
    .Q(\data_array.data1[9][26] ));
 sky130_fd_sc_hd__dfxtp_2 _12475_ (.CLK(clk),
    .D(_01169_),
    .Q(\data_array.data1[9][27] ));
 sky130_fd_sc_hd__dfxtp_2 _12476_ (.CLK(clk),
    .D(_01170_),
    .Q(\data_array.data1[9][28] ));
 sky130_fd_sc_hd__dfxtp_2 _12477_ (.CLK(clk),
    .D(_01171_),
    .Q(\data_array.data1[9][29] ));
 sky130_fd_sc_hd__dfxtp_2 _12478_ (.CLK(clk),
    .D(_01172_),
    .Q(\data_array.data1[9][30] ));
 sky130_fd_sc_hd__dfxtp_2 _12479_ (.CLK(clk),
    .D(_01173_),
    .Q(\data_array.data1[9][31] ));
 sky130_fd_sc_hd__dfxtp_2 _12480_ (.CLK(clk),
    .D(_01174_),
    .Q(\data_array.data1[9][32] ));
 sky130_fd_sc_hd__dfxtp_2 _12481_ (.CLK(clk),
    .D(_01175_),
    .Q(\data_array.data1[9][33] ));
 sky130_fd_sc_hd__dfxtp_2 _12482_ (.CLK(clk),
    .D(_01176_),
    .Q(\data_array.data1[9][34] ));
 sky130_fd_sc_hd__dfxtp_2 _12483_ (.CLK(clk),
    .D(_01177_),
    .Q(\data_array.data1[9][35] ));
 sky130_fd_sc_hd__dfxtp_2 _12484_ (.CLK(clk),
    .D(_01178_),
    .Q(\data_array.data1[9][36] ));
 sky130_fd_sc_hd__dfxtp_2 _12485_ (.CLK(clk),
    .D(_01179_),
    .Q(\data_array.data1[9][37] ));
 sky130_fd_sc_hd__dfxtp_2 _12486_ (.CLK(clk),
    .D(_01180_),
    .Q(\data_array.data1[9][38] ));
 sky130_fd_sc_hd__dfxtp_2 _12487_ (.CLK(clk),
    .D(_01181_),
    .Q(\data_array.data1[9][39] ));
 sky130_fd_sc_hd__dfxtp_2 _12488_ (.CLK(clk),
    .D(_01182_),
    .Q(\data_array.data1[9][40] ));
 sky130_fd_sc_hd__dfxtp_2 _12489_ (.CLK(clk),
    .D(_01183_),
    .Q(\data_array.data1[9][41] ));
 sky130_fd_sc_hd__dfxtp_2 _12490_ (.CLK(clk),
    .D(_01184_),
    .Q(\data_array.data1[9][42] ));
 sky130_fd_sc_hd__dfxtp_2 _12491_ (.CLK(clk),
    .D(_01185_),
    .Q(\data_array.data1[9][43] ));
 sky130_fd_sc_hd__dfxtp_2 _12492_ (.CLK(clk),
    .D(_01186_),
    .Q(\data_array.data1[9][44] ));
 sky130_fd_sc_hd__dfxtp_2 _12493_ (.CLK(clk),
    .D(_01187_),
    .Q(\data_array.data1[9][45] ));
 sky130_fd_sc_hd__dfxtp_2 _12494_ (.CLK(clk),
    .D(_01188_),
    .Q(\data_array.data1[9][46] ));
 sky130_fd_sc_hd__dfxtp_2 _12495_ (.CLK(clk),
    .D(_01189_),
    .Q(\data_array.data1[9][47] ));
 sky130_fd_sc_hd__dfxtp_2 _12496_ (.CLK(clk),
    .D(_01190_),
    .Q(\data_array.data1[9][48] ));
 sky130_fd_sc_hd__dfxtp_2 _12497_ (.CLK(clk),
    .D(_01191_),
    .Q(\data_array.data1[9][49] ));
 sky130_fd_sc_hd__dfxtp_2 _12498_ (.CLK(clk),
    .D(_01192_),
    .Q(\data_array.data1[9][50] ));
 sky130_fd_sc_hd__dfxtp_2 _12499_ (.CLK(clk),
    .D(_01193_),
    .Q(\data_array.data1[9][51] ));
 sky130_fd_sc_hd__dfxtp_2 _12500_ (.CLK(clk),
    .D(_01194_),
    .Q(\data_array.data1[9][52] ));
 sky130_fd_sc_hd__dfxtp_2 _12501_ (.CLK(clk),
    .D(_01195_),
    .Q(\data_array.data1[9][53] ));
 sky130_fd_sc_hd__dfxtp_2 _12502_ (.CLK(clk),
    .D(_01196_),
    .Q(\data_array.data1[9][54] ));
 sky130_fd_sc_hd__dfxtp_2 _12503_ (.CLK(clk),
    .D(_01197_),
    .Q(\data_array.data1[9][55] ));
 sky130_fd_sc_hd__dfxtp_2 _12504_ (.CLK(clk),
    .D(_01198_),
    .Q(\data_array.data1[9][56] ));
 sky130_fd_sc_hd__dfxtp_2 _12505_ (.CLK(clk),
    .D(_01199_),
    .Q(\data_array.data1[9][57] ));
 sky130_fd_sc_hd__dfxtp_2 _12506_ (.CLK(clk),
    .D(_01200_),
    .Q(\data_array.data1[9][58] ));
 sky130_fd_sc_hd__dfxtp_2 _12507_ (.CLK(clk),
    .D(_01201_),
    .Q(\data_array.data1[9][59] ));
 sky130_fd_sc_hd__dfxtp_2 _12508_ (.CLK(clk),
    .D(_01202_),
    .Q(\data_array.data1[9][60] ));
 sky130_fd_sc_hd__dfxtp_2 _12509_ (.CLK(clk),
    .D(_01203_),
    .Q(\data_array.data1[9][61] ));
 sky130_fd_sc_hd__dfxtp_2 _12510_ (.CLK(clk),
    .D(_01204_),
    .Q(\data_array.data1[9][62] ));
 sky130_fd_sc_hd__dfxtp_2 _12511_ (.CLK(clk),
    .D(_01205_),
    .Q(\data_array.data1[9][63] ));
 sky130_fd_sc_hd__dfxtp_2 _12512_ (.CLK(clk),
    .D(_01206_),
    .Q(\lru_array.lru_mem[8] ));
 sky130_fd_sc_hd__dfxtp_2 _12513_ (.CLK(clk),
    .D(_01207_),
    .Q(\lru_array.lru_mem[0] ));
 sky130_fd_sc_hd__dfxtp_2 _12514_ (.CLK(clk),
    .D(_01208_),
    .Q(\lru_array.lru_mem[15] ));
 sky130_fd_sc_hd__dfxtp_2 _12515_ (.CLK(clk),
    .D(_01209_),
    .Q(\lru_array.lru_mem[10] ));
 sky130_fd_sc_hd__dfxtp_2 _12516_ (.CLK(clk),
    .D(_01210_),
    .Q(\lru_array.lru_mem[1] ));
 sky130_fd_sc_hd__dfxtp_2 _12517_ (.CLK(clk),
    .D(_01211_),
    .Q(\lru_array.lru_mem[11] ));
 sky130_fd_sc_hd__dfxtp_2 _12518_ (.CLK(clk),
    .D(_01212_),
    .Q(\tag_array.tag1[11][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12519_ (.CLK(clk),
    .D(_01213_),
    .Q(\tag_array.tag1[11][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12520_ (.CLK(clk),
    .D(_01214_),
    .Q(\tag_array.tag1[11][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12521_ (.CLK(clk),
    .D(_01215_),
    .Q(\tag_array.tag1[11][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12522_ (.CLK(clk),
    .D(_01216_),
    .Q(\tag_array.tag1[11][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12523_ (.CLK(clk),
    .D(_01217_),
    .Q(\tag_array.tag1[11][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12524_ (.CLK(clk),
    .D(_01218_),
    .Q(\tag_array.tag1[11][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12525_ (.CLK(clk),
    .D(_01219_),
    .Q(\tag_array.tag1[11][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12526_ (.CLK(clk),
    .D(_01220_),
    .Q(\tag_array.tag1[11][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12527_ (.CLK(clk),
    .D(_01221_),
    .Q(\tag_array.tag1[11][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12528_ (.CLK(clk),
    .D(_01222_),
    .Q(\tag_array.tag1[11][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12529_ (.CLK(clk),
    .D(_01223_),
    .Q(\tag_array.tag1[11][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12530_ (.CLK(clk),
    .D(_01224_),
    .Q(\tag_array.tag1[11][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12531_ (.CLK(clk),
    .D(_01225_),
    .Q(\tag_array.tag1[11][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12532_ (.CLK(clk),
    .D(_01226_),
    .Q(\tag_array.tag1[11][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12533_ (.CLK(clk),
    .D(_01227_),
    .Q(\tag_array.tag1[11][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12534_ (.CLK(clk),
    .D(_01228_),
    .Q(\tag_array.tag1[11][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12535_ (.CLK(clk),
    .D(_01229_),
    .Q(\tag_array.tag1[11][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12536_ (.CLK(clk),
    .D(_01230_),
    .Q(\tag_array.tag1[11][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12537_ (.CLK(clk),
    .D(_01231_),
    .Q(\tag_array.tag1[11][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12538_ (.CLK(clk),
    .D(_01232_),
    .Q(\tag_array.tag1[11][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12539_ (.CLK(clk),
    .D(_01233_),
    .Q(\tag_array.tag1[11][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12540_ (.CLK(clk),
    .D(_01234_),
    .Q(\tag_array.tag1[11][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12541_ (.CLK(clk),
    .D(_01235_),
    .Q(\tag_array.tag1[11][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12542_ (.CLK(clk),
    .D(_01236_),
    .Q(\tag_array.tag1[11][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12543_ (.CLK(clk),
    .D(_01237_),
    .Q(\tag_array.tag0[11][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12544_ (.CLK(clk),
    .D(_01238_),
    .Q(\tag_array.tag0[11][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12545_ (.CLK(clk),
    .D(_01239_),
    .Q(\tag_array.tag0[11][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12546_ (.CLK(clk),
    .D(_01240_),
    .Q(\tag_array.tag0[11][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12547_ (.CLK(clk),
    .D(_01241_),
    .Q(\tag_array.tag0[11][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12548_ (.CLK(clk),
    .D(_01242_),
    .Q(\tag_array.tag0[11][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12549_ (.CLK(clk),
    .D(_01243_),
    .Q(\tag_array.tag0[11][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12550_ (.CLK(clk),
    .D(_01244_),
    .Q(\tag_array.tag0[11][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12551_ (.CLK(clk),
    .D(_01245_),
    .Q(\tag_array.tag0[11][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12552_ (.CLK(clk),
    .D(_01246_),
    .Q(\tag_array.tag0[11][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12553_ (.CLK(clk),
    .D(_01247_),
    .Q(\tag_array.tag0[11][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12554_ (.CLK(clk),
    .D(_01248_),
    .Q(\tag_array.tag0[11][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12555_ (.CLK(clk),
    .D(_01249_),
    .Q(\tag_array.tag0[11][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12556_ (.CLK(clk),
    .D(_01250_),
    .Q(\tag_array.tag0[11][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12557_ (.CLK(clk),
    .D(_01251_),
    .Q(\tag_array.tag0[11][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12558_ (.CLK(clk),
    .D(_01252_),
    .Q(\tag_array.tag0[11][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12559_ (.CLK(clk),
    .D(_01253_),
    .Q(\tag_array.tag0[11][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12560_ (.CLK(clk),
    .D(_01254_),
    .Q(\tag_array.tag0[11][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12561_ (.CLK(clk),
    .D(_01255_),
    .Q(\tag_array.tag0[11][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12562_ (.CLK(clk),
    .D(_01256_),
    .Q(\tag_array.tag0[11][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12563_ (.CLK(clk),
    .D(_01257_),
    .Q(\tag_array.tag0[11][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12564_ (.CLK(clk),
    .D(_01258_),
    .Q(\tag_array.tag0[11][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12565_ (.CLK(clk),
    .D(_01259_),
    .Q(\tag_array.tag0[11][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12566_ (.CLK(clk),
    .D(_01260_),
    .Q(\tag_array.tag0[11][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12567_ (.CLK(clk),
    .D(_01261_),
    .Q(\tag_array.tag0[11][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12568_ (.CLK(clk),
    .D(_01262_),
    .Q(\tag_array.tag0[10][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12569_ (.CLK(clk),
    .D(_01263_),
    .Q(\tag_array.tag0[10][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12570_ (.CLK(clk),
    .D(_01264_),
    .Q(\tag_array.tag0[10][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12571_ (.CLK(clk),
    .D(_01265_),
    .Q(\tag_array.tag0[10][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12572_ (.CLK(clk),
    .D(_01266_),
    .Q(\tag_array.tag0[10][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12573_ (.CLK(clk),
    .D(_01267_),
    .Q(\tag_array.tag0[10][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12574_ (.CLK(clk),
    .D(_01268_),
    .Q(\tag_array.tag0[10][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12575_ (.CLK(clk),
    .D(_01269_),
    .Q(\tag_array.tag0[10][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12576_ (.CLK(clk),
    .D(_01270_),
    .Q(\tag_array.tag0[10][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12577_ (.CLK(clk),
    .D(_01271_),
    .Q(\tag_array.tag0[10][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12578_ (.CLK(clk),
    .D(_01272_),
    .Q(\tag_array.tag0[10][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12579_ (.CLK(clk),
    .D(_01273_),
    .Q(\tag_array.tag0[10][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12580_ (.CLK(clk),
    .D(_01274_),
    .Q(\tag_array.tag0[10][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12581_ (.CLK(clk),
    .D(_01275_),
    .Q(\tag_array.tag0[10][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12582_ (.CLK(clk),
    .D(_01276_),
    .Q(\tag_array.tag0[10][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12583_ (.CLK(clk),
    .D(_01277_),
    .Q(\tag_array.tag0[10][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12584_ (.CLK(clk),
    .D(_01278_),
    .Q(\tag_array.tag0[10][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12585_ (.CLK(clk),
    .D(_01279_),
    .Q(\tag_array.tag0[10][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12586_ (.CLK(clk),
    .D(_01280_),
    .Q(\tag_array.tag0[10][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12587_ (.CLK(clk),
    .D(_01281_),
    .Q(\tag_array.tag0[10][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12588_ (.CLK(clk),
    .D(_01282_),
    .Q(\tag_array.tag0[10][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12589_ (.CLK(clk),
    .D(_01283_),
    .Q(\tag_array.tag0[10][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12590_ (.CLK(clk),
    .D(_01284_),
    .Q(\tag_array.tag0[10][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12591_ (.CLK(clk),
    .D(_01285_),
    .Q(\tag_array.tag0[10][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12592_ (.CLK(clk),
    .D(_01286_),
    .Q(\tag_array.tag0[10][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12593_ (.CLK(clk),
    .D(_01287_),
    .Q(\tag_array.tag0[0][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12594_ (.CLK(clk),
    .D(_01288_),
    .Q(\tag_array.tag0[0][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12595_ (.CLK(clk),
    .D(_01289_),
    .Q(\tag_array.tag0[0][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12596_ (.CLK(clk),
    .D(_01290_),
    .Q(\tag_array.tag0[0][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12597_ (.CLK(clk),
    .D(_01291_),
    .Q(\tag_array.tag0[0][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12598_ (.CLK(clk),
    .D(_01292_),
    .Q(\tag_array.tag0[0][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12599_ (.CLK(clk),
    .D(_01293_),
    .Q(\tag_array.tag0[0][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12600_ (.CLK(clk),
    .D(_01294_),
    .Q(\tag_array.tag0[0][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12601_ (.CLK(clk),
    .D(_01295_),
    .Q(\tag_array.tag0[0][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12602_ (.CLK(clk),
    .D(_01296_),
    .Q(\tag_array.tag0[0][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12603_ (.CLK(clk),
    .D(_01297_),
    .Q(\tag_array.tag0[0][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12604_ (.CLK(clk),
    .D(_01298_),
    .Q(\tag_array.tag0[0][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12605_ (.CLK(clk),
    .D(_01299_),
    .Q(\tag_array.tag0[0][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12606_ (.CLK(clk),
    .D(_01300_),
    .Q(\tag_array.tag0[0][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12607_ (.CLK(clk),
    .D(_01301_),
    .Q(\tag_array.tag0[0][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12608_ (.CLK(clk),
    .D(_01302_),
    .Q(\tag_array.tag0[0][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12609_ (.CLK(clk),
    .D(_01303_),
    .Q(\tag_array.tag0[0][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12610_ (.CLK(clk),
    .D(_01304_),
    .Q(\tag_array.tag0[0][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12611_ (.CLK(clk),
    .D(_01305_),
    .Q(\tag_array.tag0[0][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12612_ (.CLK(clk),
    .D(_01306_),
    .Q(\tag_array.tag0[0][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12613_ (.CLK(clk),
    .D(_01307_),
    .Q(\tag_array.tag0[0][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12614_ (.CLK(clk),
    .D(_01308_),
    .Q(\tag_array.tag0[0][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12615_ (.CLK(clk),
    .D(_01309_),
    .Q(\tag_array.tag0[0][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12616_ (.CLK(clk),
    .D(_01310_),
    .Q(\tag_array.tag0[0][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12617_ (.CLK(clk),
    .D(_01311_),
    .Q(\tag_array.tag0[0][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12618_ (.CLK(clk),
    .D(_01312_),
    .Q(\data_array.data0[15][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12619_ (.CLK(clk),
    .D(_01313_),
    .Q(\data_array.data0[15][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12620_ (.CLK(clk),
    .D(_01314_),
    .Q(\data_array.data0[15][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12621_ (.CLK(clk),
    .D(_01315_),
    .Q(\data_array.data0[15][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12622_ (.CLK(clk),
    .D(_01316_),
    .Q(\data_array.data0[15][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12623_ (.CLK(clk),
    .D(_01317_),
    .Q(\data_array.data0[15][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12624_ (.CLK(clk),
    .D(_01318_),
    .Q(\data_array.data0[15][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12625_ (.CLK(clk),
    .D(_01319_),
    .Q(\data_array.data0[15][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12626_ (.CLK(clk),
    .D(_01320_),
    .Q(\data_array.data0[15][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12627_ (.CLK(clk),
    .D(_01321_),
    .Q(\data_array.data0[15][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12628_ (.CLK(clk),
    .D(_01322_),
    .Q(\data_array.data0[15][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12629_ (.CLK(clk),
    .D(_01323_),
    .Q(\data_array.data0[15][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12630_ (.CLK(clk),
    .D(_01324_),
    .Q(\data_array.data0[15][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12631_ (.CLK(clk),
    .D(_01325_),
    .Q(\data_array.data0[15][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12632_ (.CLK(clk),
    .D(_01326_),
    .Q(\data_array.data0[15][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12633_ (.CLK(clk),
    .D(_01327_),
    .Q(\data_array.data0[15][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12634_ (.CLK(clk),
    .D(_01328_),
    .Q(\data_array.data0[15][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12635_ (.CLK(clk),
    .D(_01329_),
    .Q(\data_array.data0[15][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12636_ (.CLK(clk),
    .D(_01330_),
    .Q(\data_array.data0[15][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12637_ (.CLK(clk),
    .D(_01331_),
    .Q(\data_array.data0[15][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12638_ (.CLK(clk),
    .D(_01332_),
    .Q(\data_array.data0[15][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12639_ (.CLK(clk),
    .D(_01333_),
    .Q(\data_array.data0[15][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12640_ (.CLK(clk),
    .D(_01334_),
    .Q(\data_array.data0[15][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12641_ (.CLK(clk),
    .D(_01335_),
    .Q(\data_array.data0[15][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12642_ (.CLK(clk),
    .D(_01336_),
    .Q(\data_array.data0[15][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12643_ (.CLK(clk),
    .D(_01337_),
    .Q(\data_array.data0[15][25] ));
 sky130_fd_sc_hd__dfxtp_2 _12644_ (.CLK(clk),
    .D(_01338_),
    .Q(\data_array.data0[15][26] ));
 sky130_fd_sc_hd__dfxtp_2 _12645_ (.CLK(clk),
    .D(_01339_),
    .Q(\data_array.data0[15][27] ));
 sky130_fd_sc_hd__dfxtp_2 _12646_ (.CLK(clk),
    .D(_01340_),
    .Q(\data_array.data0[15][28] ));
 sky130_fd_sc_hd__dfxtp_2 _12647_ (.CLK(clk),
    .D(_01341_),
    .Q(\data_array.data0[15][29] ));
 sky130_fd_sc_hd__dfxtp_2 _12648_ (.CLK(clk),
    .D(_01342_),
    .Q(\data_array.data0[15][30] ));
 sky130_fd_sc_hd__dfxtp_2 _12649_ (.CLK(clk),
    .D(_01343_),
    .Q(\data_array.data0[15][31] ));
 sky130_fd_sc_hd__dfxtp_2 _12650_ (.CLK(clk),
    .D(_01344_),
    .Q(\data_array.data0[15][32] ));
 sky130_fd_sc_hd__dfxtp_2 _12651_ (.CLK(clk),
    .D(_01345_),
    .Q(\data_array.data0[15][33] ));
 sky130_fd_sc_hd__dfxtp_2 _12652_ (.CLK(clk),
    .D(_01346_),
    .Q(\data_array.data0[15][34] ));
 sky130_fd_sc_hd__dfxtp_2 _12653_ (.CLK(clk),
    .D(_01347_),
    .Q(\data_array.data0[15][35] ));
 sky130_fd_sc_hd__dfxtp_2 _12654_ (.CLK(clk),
    .D(_01348_),
    .Q(\data_array.data0[15][36] ));
 sky130_fd_sc_hd__dfxtp_2 _12655_ (.CLK(clk),
    .D(_01349_),
    .Q(\data_array.data0[15][37] ));
 sky130_fd_sc_hd__dfxtp_2 _12656_ (.CLK(clk),
    .D(_01350_),
    .Q(\data_array.data0[15][38] ));
 sky130_fd_sc_hd__dfxtp_2 _12657_ (.CLK(clk),
    .D(_01351_),
    .Q(\data_array.data0[15][39] ));
 sky130_fd_sc_hd__dfxtp_2 _12658_ (.CLK(clk),
    .D(_01352_),
    .Q(\data_array.data0[15][40] ));
 sky130_fd_sc_hd__dfxtp_2 _12659_ (.CLK(clk),
    .D(_01353_),
    .Q(\data_array.data0[15][41] ));
 sky130_fd_sc_hd__dfxtp_2 _12660_ (.CLK(clk),
    .D(_01354_),
    .Q(\data_array.data0[15][42] ));
 sky130_fd_sc_hd__dfxtp_2 _12661_ (.CLK(clk),
    .D(_01355_),
    .Q(\data_array.data0[15][43] ));
 sky130_fd_sc_hd__dfxtp_2 _12662_ (.CLK(clk),
    .D(_01356_),
    .Q(\data_array.data0[15][44] ));
 sky130_fd_sc_hd__dfxtp_2 _12663_ (.CLK(clk),
    .D(_01357_),
    .Q(\data_array.data0[15][45] ));
 sky130_fd_sc_hd__dfxtp_2 _12664_ (.CLK(clk),
    .D(_01358_),
    .Q(\data_array.data0[15][46] ));
 sky130_fd_sc_hd__dfxtp_2 _12665_ (.CLK(clk),
    .D(_01359_),
    .Q(\data_array.data0[15][47] ));
 sky130_fd_sc_hd__dfxtp_2 _12666_ (.CLK(clk),
    .D(_01360_),
    .Q(\data_array.data0[15][48] ));
 sky130_fd_sc_hd__dfxtp_2 _12667_ (.CLK(clk),
    .D(_01361_),
    .Q(\data_array.data0[15][49] ));
 sky130_fd_sc_hd__dfxtp_2 _12668_ (.CLK(clk),
    .D(_01362_),
    .Q(\data_array.data0[15][50] ));
 sky130_fd_sc_hd__dfxtp_2 _12669_ (.CLK(clk),
    .D(_01363_),
    .Q(\data_array.data0[15][51] ));
 sky130_fd_sc_hd__dfxtp_2 _12670_ (.CLK(clk),
    .D(_01364_),
    .Q(\data_array.data0[15][52] ));
 sky130_fd_sc_hd__dfxtp_2 _12671_ (.CLK(clk),
    .D(_01365_),
    .Q(\data_array.data0[15][53] ));
 sky130_fd_sc_hd__dfxtp_2 _12672_ (.CLK(clk),
    .D(_01366_),
    .Q(\data_array.data0[15][54] ));
 sky130_fd_sc_hd__dfxtp_2 _12673_ (.CLK(clk),
    .D(_01367_),
    .Q(\data_array.data0[15][55] ));
 sky130_fd_sc_hd__dfxtp_2 _12674_ (.CLK(clk),
    .D(_01368_),
    .Q(\data_array.data0[15][56] ));
 sky130_fd_sc_hd__dfxtp_2 _12675_ (.CLK(clk),
    .D(_01369_),
    .Q(\data_array.data0[15][57] ));
 sky130_fd_sc_hd__dfxtp_2 _12676_ (.CLK(clk),
    .D(_01370_),
    .Q(\data_array.data0[15][58] ));
 sky130_fd_sc_hd__dfxtp_2 _12677_ (.CLK(clk),
    .D(_01371_),
    .Q(\data_array.data0[15][59] ));
 sky130_fd_sc_hd__dfxtp_2 _12678_ (.CLK(clk),
    .D(_01372_),
    .Q(\data_array.data0[15][60] ));
 sky130_fd_sc_hd__dfxtp_2 _12679_ (.CLK(clk),
    .D(_01373_),
    .Q(\data_array.data0[15][61] ));
 sky130_fd_sc_hd__dfxtp_2 _12680_ (.CLK(clk),
    .D(_01374_),
    .Q(\data_array.data0[15][62] ));
 sky130_fd_sc_hd__dfxtp_2 _12681_ (.CLK(clk),
    .D(_01375_),
    .Q(\data_array.data0[15][63] ));
 sky130_fd_sc_hd__dfxtp_2 _12682_ (.CLK(clk),
    .D(_01376_),
    .Q(\tag_array.tag0[8][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12683_ (.CLK(clk),
    .D(_01377_),
    .Q(\tag_array.tag0[8][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12684_ (.CLK(clk),
    .D(_01378_),
    .Q(\tag_array.tag0[8][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12685_ (.CLK(clk),
    .D(_01379_),
    .Q(\tag_array.tag0[8][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12686_ (.CLK(clk),
    .D(_01380_),
    .Q(\tag_array.tag0[8][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12687_ (.CLK(clk),
    .D(_01381_),
    .Q(\tag_array.tag0[8][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12688_ (.CLK(clk),
    .D(_01382_),
    .Q(\tag_array.tag0[8][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12689_ (.CLK(clk),
    .D(_01383_),
    .Q(\tag_array.tag0[8][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12690_ (.CLK(clk),
    .D(_01384_),
    .Q(\tag_array.tag0[8][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12691_ (.CLK(clk),
    .D(_01385_),
    .Q(\tag_array.tag0[8][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12692_ (.CLK(clk),
    .D(_01386_),
    .Q(\tag_array.tag0[8][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12693_ (.CLK(clk),
    .D(_01387_),
    .Q(\tag_array.tag0[8][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12694_ (.CLK(clk),
    .D(_01388_),
    .Q(\tag_array.tag0[8][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12695_ (.CLK(clk),
    .D(_01389_),
    .Q(\tag_array.tag0[8][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12696_ (.CLK(clk),
    .D(_01390_),
    .Q(\tag_array.tag0[8][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12697_ (.CLK(clk),
    .D(_01391_),
    .Q(\tag_array.tag0[8][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12698_ (.CLK(clk),
    .D(_01392_),
    .Q(\tag_array.tag0[8][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12699_ (.CLK(clk),
    .D(_01393_),
    .Q(\tag_array.tag0[8][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12700_ (.CLK(clk),
    .D(_01394_),
    .Q(\tag_array.tag0[8][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12701_ (.CLK(clk),
    .D(_01395_),
    .Q(\tag_array.tag0[8][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12702_ (.CLK(clk),
    .D(_01396_),
    .Q(\tag_array.tag0[8][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12703_ (.CLK(clk),
    .D(_01397_),
    .Q(\tag_array.tag0[8][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12704_ (.CLK(clk),
    .D(_01398_),
    .Q(\tag_array.tag0[8][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12705_ (.CLK(clk),
    .D(_01399_),
    .Q(\tag_array.tag0[8][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12706_ (.CLK(clk),
    .D(_01400_),
    .Q(\tag_array.tag0[8][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12707_ (.CLK(clk),
    .D(_01401_),
    .Q(\tag_array.tag0[7][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12708_ (.CLK(clk),
    .D(_01402_),
    .Q(\tag_array.tag0[7][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12709_ (.CLK(clk),
    .D(_01403_),
    .Q(\tag_array.tag0[7][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12710_ (.CLK(clk),
    .D(_01404_),
    .Q(\tag_array.tag0[7][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12711_ (.CLK(clk),
    .D(_01405_),
    .Q(\tag_array.tag0[7][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12712_ (.CLK(clk),
    .D(_01406_),
    .Q(\tag_array.tag0[7][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12713_ (.CLK(clk),
    .D(_01407_),
    .Q(\tag_array.tag0[7][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12714_ (.CLK(clk),
    .D(_01408_),
    .Q(\tag_array.tag0[7][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12715_ (.CLK(clk),
    .D(_01409_),
    .Q(\tag_array.tag0[7][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12716_ (.CLK(clk),
    .D(_01410_),
    .Q(\tag_array.tag0[7][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12717_ (.CLK(clk),
    .D(_01411_),
    .Q(\tag_array.tag0[7][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12718_ (.CLK(clk),
    .D(_01412_),
    .Q(\tag_array.tag0[7][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12719_ (.CLK(clk),
    .D(_01413_),
    .Q(\tag_array.tag0[7][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12720_ (.CLK(clk),
    .D(_01414_),
    .Q(\tag_array.tag0[7][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12721_ (.CLK(clk),
    .D(_01415_),
    .Q(\tag_array.tag0[7][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12722_ (.CLK(clk),
    .D(_01416_),
    .Q(\tag_array.tag0[7][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12723_ (.CLK(clk),
    .D(_01417_),
    .Q(\tag_array.tag0[7][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12724_ (.CLK(clk),
    .D(_01418_),
    .Q(\tag_array.tag0[7][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12725_ (.CLK(clk),
    .D(_01419_),
    .Q(\tag_array.tag0[7][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12726_ (.CLK(clk),
    .D(_01420_),
    .Q(\tag_array.tag0[7][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12727_ (.CLK(clk),
    .D(_01421_),
    .Q(\tag_array.tag0[7][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12728_ (.CLK(clk),
    .D(_01422_),
    .Q(\tag_array.tag0[7][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12729_ (.CLK(clk),
    .D(_01423_),
    .Q(\tag_array.tag0[7][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12730_ (.CLK(clk),
    .D(_01424_),
    .Q(\tag_array.tag0[7][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12731_ (.CLK(clk),
    .D(_01425_),
    .Q(\tag_array.tag0[7][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12732_ (.CLK(clk),
    .D(_01426_),
    .Q(\tag_array.tag0[5][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12733_ (.CLK(clk),
    .D(_01427_),
    .Q(\tag_array.tag0[5][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12734_ (.CLK(clk),
    .D(_01428_),
    .Q(\tag_array.tag0[5][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12735_ (.CLK(clk),
    .D(_01429_),
    .Q(\tag_array.tag0[5][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12736_ (.CLK(clk),
    .D(_01430_),
    .Q(\tag_array.tag0[5][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12737_ (.CLK(clk),
    .D(_01431_),
    .Q(\tag_array.tag0[5][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12738_ (.CLK(clk),
    .D(_01432_),
    .Q(\tag_array.tag0[5][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12739_ (.CLK(clk),
    .D(_01433_),
    .Q(\tag_array.tag0[5][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12740_ (.CLK(clk),
    .D(_01434_),
    .Q(\tag_array.tag0[5][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12741_ (.CLK(clk),
    .D(_01435_),
    .Q(\tag_array.tag0[5][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12742_ (.CLK(clk),
    .D(_01436_),
    .Q(\tag_array.tag0[5][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12743_ (.CLK(clk),
    .D(_01437_),
    .Q(\tag_array.tag0[5][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12744_ (.CLK(clk),
    .D(_01438_),
    .Q(\tag_array.tag0[5][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12745_ (.CLK(clk),
    .D(_01439_),
    .Q(\tag_array.tag0[5][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12746_ (.CLK(clk),
    .D(_01440_),
    .Q(\tag_array.tag0[5][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12747_ (.CLK(clk),
    .D(_01441_),
    .Q(\tag_array.tag0[5][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12748_ (.CLK(clk),
    .D(_01442_),
    .Q(\tag_array.tag0[5][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12749_ (.CLK(clk),
    .D(_01443_),
    .Q(\tag_array.tag0[5][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12750_ (.CLK(clk),
    .D(_01444_),
    .Q(\tag_array.tag0[5][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12751_ (.CLK(clk),
    .D(_01445_),
    .Q(\tag_array.tag0[5][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12752_ (.CLK(clk),
    .D(_01446_),
    .Q(\tag_array.tag0[5][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12753_ (.CLK(clk),
    .D(_01447_),
    .Q(\tag_array.tag0[5][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12754_ (.CLK(clk),
    .D(_01448_),
    .Q(\tag_array.tag0[5][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12755_ (.CLK(clk),
    .D(_01449_),
    .Q(\tag_array.tag0[5][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12756_ (.CLK(clk),
    .D(_01450_),
    .Q(\tag_array.tag0[5][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12757_ (.CLK(clk),
    .D(_01451_),
    .Q(\tag_array.tag0[6][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12758_ (.CLK(clk),
    .D(_01452_),
    .Q(\tag_array.tag0[6][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12759_ (.CLK(clk),
    .D(_01453_),
    .Q(\tag_array.tag0[6][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12760_ (.CLK(clk),
    .D(_01454_),
    .Q(\tag_array.tag0[6][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12761_ (.CLK(clk),
    .D(_01455_),
    .Q(\tag_array.tag0[6][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12762_ (.CLK(clk),
    .D(_01456_),
    .Q(\tag_array.tag0[6][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12763_ (.CLK(clk),
    .D(_01457_),
    .Q(\tag_array.tag0[6][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12764_ (.CLK(clk),
    .D(_01458_),
    .Q(\tag_array.tag0[6][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12765_ (.CLK(clk),
    .D(_01459_),
    .Q(\tag_array.tag0[6][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12766_ (.CLK(clk),
    .D(_01460_),
    .Q(\tag_array.tag0[6][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12767_ (.CLK(clk),
    .D(_01461_),
    .Q(\tag_array.tag0[6][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12768_ (.CLK(clk),
    .D(_01462_),
    .Q(\tag_array.tag0[6][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12769_ (.CLK(clk),
    .D(_01463_),
    .Q(\tag_array.tag0[6][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12770_ (.CLK(clk),
    .D(_01464_),
    .Q(\tag_array.tag0[6][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12771_ (.CLK(clk),
    .D(_01465_),
    .Q(\tag_array.tag0[6][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12772_ (.CLK(clk),
    .D(_01466_),
    .Q(\tag_array.tag0[6][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12773_ (.CLK(clk),
    .D(_01467_),
    .Q(\tag_array.tag0[6][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12774_ (.CLK(clk),
    .D(_01468_),
    .Q(\tag_array.tag0[6][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12775_ (.CLK(clk),
    .D(_01469_),
    .Q(\tag_array.tag0[6][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12776_ (.CLK(clk),
    .D(_01470_),
    .Q(\tag_array.tag0[6][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12777_ (.CLK(clk),
    .D(_01471_),
    .Q(\tag_array.tag0[6][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12778_ (.CLK(clk),
    .D(_01472_),
    .Q(\tag_array.tag0[6][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12779_ (.CLK(clk),
    .D(_01473_),
    .Q(\tag_array.tag0[6][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12780_ (.CLK(clk),
    .D(_01474_),
    .Q(\tag_array.tag0[6][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12781_ (.CLK(clk),
    .D(_01475_),
    .Q(\tag_array.tag0[6][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12782_ (.CLK(clk),
    .D(_01476_),
    .Q(\tag_array.tag1[10][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12783_ (.CLK(clk),
    .D(_01477_),
    .Q(\tag_array.tag1[10][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12784_ (.CLK(clk),
    .D(_01478_),
    .Q(\tag_array.tag1[10][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12785_ (.CLK(clk),
    .D(_01479_),
    .Q(\tag_array.tag1[10][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12786_ (.CLK(clk),
    .D(_01480_),
    .Q(\tag_array.tag1[10][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12787_ (.CLK(clk),
    .D(_01481_),
    .Q(\tag_array.tag1[10][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12788_ (.CLK(clk),
    .D(_01482_),
    .Q(\tag_array.tag1[10][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12789_ (.CLK(clk),
    .D(_01483_),
    .Q(\tag_array.tag1[10][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12790_ (.CLK(clk),
    .D(_01484_),
    .Q(\tag_array.tag1[10][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12791_ (.CLK(clk),
    .D(_01485_),
    .Q(\tag_array.tag1[10][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12792_ (.CLK(clk),
    .D(_01486_),
    .Q(\tag_array.tag1[10][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12793_ (.CLK(clk),
    .D(_01487_),
    .Q(\tag_array.tag1[10][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12794_ (.CLK(clk),
    .D(_01488_),
    .Q(\tag_array.tag1[10][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12795_ (.CLK(clk),
    .D(_01489_),
    .Q(\tag_array.tag1[10][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12796_ (.CLK(clk),
    .D(_01490_),
    .Q(\tag_array.tag1[10][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12797_ (.CLK(clk),
    .D(_01491_),
    .Q(\tag_array.tag1[10][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12798_ (.CLK(clk),
    .D(_01492_),
    .Q(\tag_array.tag1[10][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12799_ (.CLK(clk),
    .D(_01493_),
    .Q(\tag_array.tag1[10][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12800_ (.CLK(clk),
    .D(_01494_),
    .Q(\tag_array.tag1[10][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12801_ (.CLK(clk),
    .D(_01495_),
    .Q(\tag_array.tag1[10][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12802_ (.CLK(clk),
    .D(_01496_),
    .Q(\tag_array.tag1[10][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12803_ (.CLK(clk),
    .D(_01497_),
    .Q(\tag_array.tag1[10][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12804_ (.CLK(clk),
    .D(_01498_),
    .Q(\tag_array.tag1[10][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12805_ (.CLK(clk),
    .D(_01499_),
    .Q(\tag_array.tag1[10][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12806_ (.CLK(clk),
    .D(_01500_),
    .Q(\tag_array.tag1[10][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12807_ (.CLK(clk),
    .D(_01501_),
    .Q(\tag_array.tag1[0][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12808_ (.CLK(clk),
    .D(_01502_),
    .Q(\tag_array.tag1[0][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12809_ (.CLK(clk),
    .D(_01503_),
    .Q(\tag_array.tag1[0][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12810_ (.CLK(clk),
    .D(_01504_),
    .Q(\tag_array.tag1[0][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12811_ (.CLK(clk),
    .D(_01505_),
    .Q(\tag_array.tag1[0][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12812_ (.CLK(clk),
    .D(_01506_),
    .Q(\tag_array.tag1[0][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12813_ (.CLK(clk),
    .D(_01507_),
    .Q(\tag_array.tag1[0][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12814_ (.CLK(clk),
    .D(_01508_),
    .Q(\tag_array.tag1[0][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12815_ (.CLK(clk),
    .D(_01509_),
    .Q(\tag_array.tag1[0][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12816_ (.CLK(clk),
    .D(_01510_),
    .Q(\tag_array.tag1[0][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12817_ (.CLK(clk),
    .D(_01511_),
    .Q(\tag_array.tag1[0][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12818_ (.CLK(clk),
    .D(_01512_),
    .Q(\tag_array.tag1[0][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12819_ (.CLK(clk),
    .D(_01513_),
    .Q(\tag_array.tag1[0][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12820_ (.CLK(clk),
    .D(_01514_),
    .Q(\tag_array.tag1[0][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12821_ (.CLK(clk),
    .D(_01515_),
    .Q(\tag_array.tag1[0][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12822_ (.CLK(clk),
    .D(_01516_),
    .Q(\tag_array.tag1[0][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12823_ (.CLK(clk),
    .D(_01517_),
    .Q(\tag_array.tag1[0][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12824_ (.CLK(clk),
    .D(_01518_),
    .Q(\tag_array.tag1[0][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12825_ (.CLK(clk),
    .D(_01519_),
    .Q(\tag_array.tag1[0][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12826_ (.CLK(clk),
    .D(_01520_),
    .Q(\tag_array.tag1[0][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12827_ (.CLK(clk),
    .D(_01521_),
    .Q(\tag_array.tag1[0][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12828_ (.CLK(clk),
    .D(_01522_),
    .Q(\tag_array.tag1[0][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12829_ (.CLK(clk),
    .D(_01523_),
    .Q(\tag_array.tag1[0][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12830_ (.CLK(clk),
    .D(_01524_),
    .Q(\tag_array.tag1[0][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12831_ (.CLK(clk),
    .D(_01525_),
    .Q(\tag_array.tag1[0][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12832_ (.CLK(clk),
    .D(_01526_),
    .Q(\data_array.data0[12][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12833_ (.CLK(clk),
    .D(_01527_),
    .Q(\data_array.data0[12][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12834_ (.CLK(clk),
    .D(_01528_),
    .Q(\data_array.data0[12][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12835_ (.CLK(clk),
    .D(_01529_),
    .Q(\data_array.data0[12][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12836_ (.CLK(clk),
    .D(_01530_),
    .Q(\data_array.data0[12][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12837_ (.CLK(clk),
    .D(_01531_),
    .Q(\data_array.data0[12][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12838_ (.CLK(clk),
    .D(_01532_),
    .Q(\data_array.data0[12][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12839_ (.CLK(clk),
    .D(_01533_),
    .Q(\data_array.data0[12][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12840_ (.CLK(clk),
    .D(_01534_),
    .Q(\data_array.data0[12][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12841_ (.CLK(clk),
    .D(_01535_),
    .Q(\data_array.data0[12][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12842_ (.CLK(clk),
    .D(_01536_),
    .Q(\data_array.data0[12][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12843_ (.CLK(clk),
    .D(_01537_),
    .Q(\data_array.data0[12][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12844_ (.CLK(clk),
    .D(_01538_),
    .Q(\data_array.data0[12][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12845_ (.CLK(clk),
    .D(_01539_),
    .Q(\data_array.data0[12][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12846_ (.CLK(clk),
    .D(_01540_),
    .Q(\data_array.data0[12][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12847_ (.CLK(clk),
    .D(_01541_),
    .Q(\data_array.data0[12][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12848_ (.CLK(clk),
    .D(_01542_),
    .Q(\data_array.data0[12][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12849_ (.CLK(clk),
    .D(_01543_),
    .Q(\data_array.data0[12][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12850_ (.CLK(clk),
    .D(_01544_),
    .Q(\data_array.data0[12][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12851_ (.CLK(clk),
    .D(_01545_),
    .Q(\data_array.data0[12][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12852_ (.CLK(clk),
    .D(_01546_),
    .Q(\data_array.data0[12][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12853_ (.CLK(clk),
    .D(_01547_),
    .Q(\data_array.data0[12][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12854_ (.CLK(clk),
    .D(_01548_),
    .Q(\data_array.data0[12][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12855_ (.CLK(clk),
    .D(_01549_),
    .Q(\data_array.data0[12][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12856_ (.CLK(clk),
    .D(_01550_),
    .Q(\data_array.data0[12][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12857_ (.CLK(clk),
    .D(_01551_),
    .Q(\data_array.data0[12][25] ));
 sky130_fd_sc_hd__dfxtp_2 _12858_ (.CLK(clk),
    .D(_01552_),
    .Q(\data_array.data0[12][26] ));
 sky130_fd_sc_hd__dfxtp_2 _12859_ (.CLK(clk),
    .D(_01553_),
    .Q(\data_array.data0[12][27] ));
 sky130_fd_sc_hd__dfxtp_2 _12860_ (.CLK(clk),
    .D(_01554_),
    .Q(\data_array.data0[12][28] ));
 sky130_fd_sc_hd__dfxtp_2 _12861_ (.CLK(clk),
    .D(_01555_),
    .Q(\data_array.data0[12][29] ));
 sky130_fd_sc_hd__dfxtp_2 _12862_ (.CLK(clk),
    .D(_01556_),
    .Q(\data_array.data0[12][30] ));
 sky130_fd_sc_hd__dfxtp_2 _12863_ (.CLK(clk),
    .D(_01557_),
    .Q(\data_array.data0[12][31] ));
 sky130_fd_sc_hd__dfxtp_2 _12864_ (.CLK(clk),
    .D(_01558_),
    .Q(\data_array.data0[12][32] ));
 sky130_fd_sc_hd__dfxtp_2 _12865_ (.CLK(clk),
    .D(_01559_),
    .Q(\data_array.data0[12][33] ));
 sky130_fd_sc_hd__dfxtp_2 _12866_ (.CLK(clk),
    .D(_01560_),
    .Q(\data_array.data0[12][34] ));
 sky130_fd_sc_hd__dfxtp_2 _12867_ (.CLK(clk),
    .D(_01561_),
    .Q(\data_array.data0[12][35] ));
 sky130_fd_sc_hd__dfxtp_2 _12868_ (.CLK(clk),
    .D(_01562_),
    .Q(\data_array.data0[12][36] ));
 sky130_fd_sc_hd__dfxtp_2 _12869_ (.CLK(clk),
    .D(_01563_),
    .Q(\data_array.data0[12][37] ));
 sky130_fd_sc_hd__dfxtp_2 _12870_ (.CLK(clk),
    .D(_01564_),
    .Q(\data_array.data0[12][38] ));
 sky130_fd_sc_hd__dfxtp_2 _12871_ (.CLK(clk),
    .D(_01565_),
    .Q(\data_array.data0[12][39] ));
 sky130_fd_sc_hd__dfxtp_2 _12872_ (.CLK(clk),
    .D(_01566_),
    .Q(\data_array.data0[12][40] ));
 sky130_fd_sc_hd__dfxtp_2 _12873_ (.CLK(clk),
    .D(_01567_),
    .Q(\data_array.data0[12][41] ));
 sky130_fd_sc_hd__dfxtp_2 _12874_ (.CLK(clk),
    .D(_01568_),
    .Q(\data_array.data0[12][42] ));
 sky130_fd_sc_hd__dfxtp_2 _12875_ (.CLK(clk),
    .D(_01569_),
    .Q(\data_array.data0[12][43] ));
 sky130_fd_sc_hd__dfxtp_2 _12876_ (.CLK(clk),
    .D(_01570_),
    .Q(\data_array.data0[12][44] ));
 sky130_fd_sc_hd__dfxtp_2 _12877_ (.CLK(clk),
    .D(_01571_),
    .Q(\data_array.data0[12][45] ));
 sky130_fd_sc_hd__dfxtp_2 _12878_ (.CLK(clk),
    .D(_01572_),
    .Q(\data_array.data0[12][46] ));
 sky130_fd_sc_hd__dfxtp_2 _12879_ (.CLK(clk),
    .D(_01573_),
    .Q(\data_array.data0[12][47] ));
 sky130_fd_sc_hd__dfxtp_2 _12880_ (.CLK(clk),
    .D(_01574_),
    .Q(\data_array.data0[12][48] ));
 sky130_fd_sc_hd__dfxtp_2 _12881_ (.CLK(clk),
    .D(_01575_),
    .Q(\data_array.data0[12][49] ));
 sky130_fd_sc_hd__dfxtp_2 _12882_ (.CLK(clk),
    .D(_01576_),
    .Q(\data_array.data0[12][50] ));
 sky130_fd_sc_hd__dfxtp_2 _12883_ (.CLK(clk),
    .D(_01577_),
    .Q(\data_array.data0[12][51] ));
 sky130_fd_sc_hd__dfxtp_2 _12884_ (.CLK(clk),
    .D(_01578_),
    .Q(\data_array.data0[12][52] ));
 sky130_fd_sc_hd__dfxtp_2 _12885_ (.CLK(clk),
    .D(_01579_),
    .Q(\data_array.data0[12][53] ));
 sky130_fd_sc_hd__dfxtp_2 _12886_ (.CLK(clk),
    .D(_01580_),
    .Q(\data_array.data0[12][54] ));
 sky130_fd_sc_hd__dfxtp_2 _12887_ (.CLK(clk),
    .D(_01581_),
    .Q(\data_array.data0[12][55] ));
 sky130_fd_sc_hd__dfxtp_2 _12888_ (.CLK(clk),
    .D(_01582_),
    .Q(\data_array.data0[12][56] ));
 sky130_fd_sc_hd__dfxtp_2 _12889_ (.CLK(clk),
    .D(_01583_),
    .Q(\data_array.data0[12][57] ));
 sky130_fd_sc_hd__dfxtp_2 _12890_ (.CLK(clk),
    .D(_01584_),
    .Q(\data_array.data0[12][58] ));
 sky130_fd_sc_hd__dfxtp_2 _12891_ (.CLK(clk),
    .D(_01585_),
    .Q(\data_array.data0[12][59] ));
 sky130_fd_sc_hd__dfxtp_2 _12892_ (.CLK(clk),
    .D(_01586_),
    .Q(\data_array.data0[12][60] ));
 sky130_fd_sc_hd__dfxtp_2 _12893_ (.CLK(clk),
    .D(_01587_),
    .Q(\data_array.data0[12][61] ));
 sky130_fd_sc_hd__dfxtp_2 _12894_ (.CLK(clk),
    .D(_01588_),
    .Q(\data_array.data0[12][62] ));
 sky130_fd_sc_hd__dfxtp_2 _12895_ (.CLK(clk),
    .D(_01589_),
    .Q(\data_array.data0[12][63] ));
 sky130_fd_sc_hd__dfxtp_2 _12896_ (.CLK(clk),
    .D(_01590_),
    .Q(\data_array.data0[13][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12897_ (.CLK(clk),
    .D(_01591_),
    .Q(\data_array.data0[13][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12898_ (.CLK(clk),
    .D(_01592_),
    .Q(\data_array.data0[13][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12899_ (.CLK(clk),
    .D(_01593_),
    .Q(\data_array.data0[13][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12900_ (.CLK(clk),
    .D(_01594_),
    .Q(\data_array.data0[13][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12901_ (.CLK(clk),
    .D(_01595_),
    .Q(\data_array.data0[13][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12902_ (.CLK(clk),
    .D(_01596_),
    .Q(\data_array.data0[13][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12903_ (.CLK(clk),
    .D(_01597_),
    .Q(\data_array.data0[13][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12904_ (.CLK(clk),
    .D(_01598_),
    .Q(\data_array.data0[13][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12905_ (.CLK(clk),
    .D(_01599_),
    .Q(\data_array.data0[13][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12906_ (.CLK(clk),
    .D(_01600_),
    .Q(\data_array.data0[13][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12907_ (.CLK(clk),
    .D(_01601_),
    .Q(\data_array.data0[13][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12908_ (.CLK(clk),
    .D(_01602_),
    .Q(\data_array.data0[13][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12909_ (.CLK(clk),
    .D(_01603_),
    .Q(\data_array.data0[13][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12910_ (.CLK(clk),
    .D(_01604_),
    .Q(\data_array.data0[13][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12911_ (.CLK(clk),
    .D(_01605_),
    .Q(\data_array.data0[13][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12912_ (.CLK(clk),
    .D(_01606_),
    .Q(\data_array.data0[13][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12913_ (.CLK(clk),
    .D(_01607_),
    .Q(\data_array.data0[13][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12914_ (.CLK(clk),
    .D(_01608_),
    .Q(\data_array.data0[13][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12915_ (.CLK(clk),
    .D(_01609_),
    .Q(\data_array.data0[13][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12916_ (.CLK(clk),
    .D(_01610_),
    .Q(\data_array.data0[13][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12917_ (.CLK(clk),
    .D(_01611_),
    .Q(\data_array.data0[13][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12918_ (.CLK(clk),
    .D(_01612_),
    .Q(\data_array.data0[13][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12919_ (.CLK(clk),
    .D(_01613_),
    .Q(\data_array.data0[13][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12920_ (.CLK(clk),
    .D(_01614_),
    .Q(\data_array.data0[13][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12921_ (.CLK(clk),
    .D(_01615_),
    .Q(\data_array.data0[13][25] ));
 sky130_fd_sc_hd__dfxtp_2 _12922_ (.CLK(clk),
    .D(_01616_),
    .Q(\data_array.data0[13][26] ));
 sky130_fd_sc_hd__dfxtp_2 _12923_ (.CLK(clk),
    .D(_01617_),
    .Q(\data_array.data0[13][27] ));
 sky130_fd_sc_hd__dfxtp_2 _12924_ (.CLK(clk),
    .D(_01618_),
    .Q(\data_array.data0[13][28] ));
 sky130_fd_sc_hd__dfxtp_2 _12925_ (.CLK(clk),
    .D(_01619_),
    .Q(\data_array.data0[13][29] ));
 sky130_fd_sc_hd__dfxtp_2 _12926_ (.CLK(clk),
    .D(_01620_),
    .Q(\data_array.data0[13][30] ));
 sky130_fd_sc_hd__dfxtp_2 _12927_ (.CLK(clk),
    .D(_01621_),
    .Q(\data_array.data0[13][31] ));
 sky130_fd_sc_hd__dfxtp_2 _12928_ (.CLK(clk),
    .D(_01622_),
    .Q(\data_array.data0[13][32] ));
 sky130_fd_sc_hd__dfxtp_2 _12929_ (.CLK(clk),
    .D(_01623_),
    .Q(\data_array.data0[13][33] ));
 sky130_fd_sc_hd__dfxtp_2 _12930_ (.CLK(clk),
    .D(_01624_),
    .Q(\data_array.data0[13][34] ));
 sky130_fd_sc_hd__dfxtp_2 _12931_ (.CLK(clk),
    .D(_01625_),
    .Q(\data_array.data0[13][35] ));
 sky130_fd_sc_hd__dfxtp_2 _12932_ (.CLK(clk),
    .D(_01626_),
    .Q(\data_array.data0[13][36] ));
 sky130_fd_sc_hd__dfxtp_2 _12933_ (.CLK(clk),
    .D(_01627_),
    .Q(\data_array.data0[13][37] ));
 sky130_fd_sc_hd__dfxtp_2 _12934_ (.CLK(clk),
    .D(_01628_),
    .Q(\data_array.data0[13][38] ));
 sky130_fd_sc_hd__dfxtp_2 _12935_ (.CLK(clk),
    .D(_01629_),
    .Q(\data_array.data0[13][39] ));
 sky130_fd_sc_hd__dfxtp_2 _12936_ (.CLK(clk),
    .D(_01630_),
    .Q(\data_array.data0[13][40] ));
 sky130_fd_sc_hd__dfxtp_2 _12937_ (.CLK(clk),
    .D(_01631_),
    .Q(\data_array.data0[13][41] ));
 sky130_fd_sc_hd__dfxtp_2 _12938_ (.CLK(clk),
    .D(_01632_),
    .Q(\data_array.data0[13][42] ));
 sky130_fd_sc_hd__dfxtp_2 _12939_ (.CLK(clk),
    .D(_01633_),
    .Q(\data_array.data0[13][43] ));
 sky130_fd_sc_hd__dfxtp_2 _12940_ (.CLK(clk),
    .D(_01634_),
    .Q(\data_array.data0[13][44] ));
 sky130_fd_sc_hd__dfxtp_2 _12941_ (.CLK(clk),
    .D(_01635_),
    .Q(\data_array.data0[13][45] ));
 sky130_fd_sc_hd__dfxtp_2 _12942_ (.CLK(clk),
    .D(_01636_),
    .Q(\data_array.data0[13][46] ));
 sky130_fd_sc_hd__dfxtp_2 _12943_ (.CLK(clk),
    .D(_01637_),
    .Q(\data_array.data0[13][47] ));
 sky130_fd_sc_hd__dfxtp_2 _12944_ (.CLK(clk),
    .D(_01638_),
    .Q(\data_array.data0[13][48] ));
 sky130_fd_sc_hd__dfxtp_2 _12945_ (.CLK(clk),
    .D(_01639_),
    .Q(\data_array.data0[13][49] ));
 sky130_fd_sc_hd__dfxtp_2 _12946_ (.CLK(clk),
    .D(_01640_),
    .Q(\data_array.data0[13][50] ));
 sky130_fd_sc_hd__dfxtp_2 _12947_ (.CLK(clk),
    .D(_01641_),
    .Q(\data_array.data0[13][51] ));
 sky130_fd_sc_hd__dfxtp_2 _12948_ (.CLK(clk),
    .D(_01642_),
    .Q(\data_array.data0[13][52] ));
 sky130_fd_sc_hd__dfxtp_2 _12949_ (.CLK(clk),
    .D(_01643_),
    .Q(\data_array.data0[13][53] ));
 sky130_fd_sc_hd__dfxtp_2 _12950_ (.CLK(clk),
    .D(_01644_),
    .Q(\data_array.data0[13][54] ));
 sky130_fd_sc_hd__dfxtp_2 _12951_ (.CLK(clk),
    .D(_01645_),
    .Q(\data_array.data0[13][55] ));
 sky130_fd_sc_hd__dfxtp_2 _12952_ (.CLK(clk),
    .D(_01646_),
    .Q(\data_array.data0[13][56] ));
 sky130_fd_sc_hd__dfxtp_2 _12953_ (.CLK(clk),
    .D(_01647_),
    .Q(\data_array.data0[13][57] ));
 sky130_fd_sc_hd__dfxtp_2 _12954_ (.CLK(clk),
    .D(_01648_),
    .Q(\data_array.data0[13][58] ));
 sky130_fd_sc_hd__dfxtp_2 _12955_ (.CLK(clk),
    .D(_01649_),
    .Q(\data_array.data0[13][59] ));
 sky130_fd_sc_hd__dfxtp_2 _12956_ (.CLK(clk),
    .D(_01650_),
    .Q(\data_array.data0[13][60] ));
 sky130_fd_sc_hd__dfxtp_2 _12957_ (.CLK(clk),
    .D(_01651_),
    .Q(\data_array.data0[13][61] ));
 sky130_fd_sc_hd__dfxtp_2 _12958_ (.CLK(clk),
    .D(_01652_),
    .Q(\data_array.data0[13][62] ));
 sky130_fd_sc_hd__dfxtp_2 _12959_ (.CLK(clk),
    .D(_01653_),
    .Q(\data_array.data0[13][63] ));
 sky130_fd_sc_hd__dfxtp_2 _12960_ (.CLK(clk),
    .D(_01654_),
    .Q(\tag_array.tag0[4][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12961_ (.CLK(clk),
    .D(_01655_),
    .Q(\tag_array.tag0[4][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12962_ (.CLK(clk),
    .D(_01656_),
    .Q(\tag_array.tag0[4][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12963_ (.CLK(clk),
    .D(_01657_),
    .Q(\tag_array.tag0[4][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12964_ (.CLK(clk),
    .D(_01658_),
    .Q(\tag_array.tag0[4][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12965_ (.CLK(clk),
    .D(_01659_),
    .Q(\tag_array.tag0[4][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12966_ (.CLK(clk),
    .D(_01660_),
    .Q(\tag_array.tag0[4][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12967_ (.CLK(clk),
    .D(_01661_),
    .Q(\tag_array.tag0[4][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12968_ (.CLK(clk),
    .D(_01662_),
    .Q(\tag_array.tag0[4][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12969_ (.CLK(clk),
    .D(_01663_),
    .Q(\tag_array.tag0[4][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12970_ (.CLK(clk),
    .D(_01664_),
    .Q(\tag_array.tag0[4][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12971_ (.CLK(clk),
    .D(_01665_),
    .Q(\tag_array.tag0[4][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12972_ (.CLK(clk),
    .D(_01666_),
    .Q(\tag_array.tag0[4][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12973_ (.CLK(clk),
    .D(_01667_),
    .Q(\tag_array.tag0[4][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12974_ (.CLK(clk),
    .D(_01668_),
    .Q(\tag_array.tag0[4][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12975_ (.CLK(clk),
    .D(_01669_),
    .Q(\tag_array.tag0[4][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12976_ (.CLK(clk),
    .D(_01670_),
    .Q(\tag_array.tag0[4][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12977_ (.CLK(clk),
    .D(_01671_),
    .Q(\tag_array.tag0[4][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12978_ (.CLK(clk),
    .D(_01672_),
    .Q(\tag_array.tag0[4][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12979_ (.CLK(clk),
    .D(_01673_),
    .Q(\tag_array.tag0[4][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12980_ (.CLK(clk),
    .D(_01674_),
    .Q(\tag_array.tag0[4][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12981_ (.CLK(clk),
    .D(_01675_),
    .Q(\tag_array.tag0[4][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12982_ (.CLK(clk),
    .D(_01676_),
    .Q(\tag_array.tag0[4][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12983_ (.CLK(clk),
    .D(_01677_),
    .Q(\tag_array.tag0[4][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12984_ (.CLK(clk),
    .D(_01678_),
    .Q(\tag_array.tag0[4][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12985_ (.CLK(clk),
    .D(_01679_),
    .Q(\data_array.data0[3][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12986_ (.CLK(clk),
    .D(_01680_),
    .Q(\data_array.data0[3][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12987_ (.CLK(clk),
    .D(_01681_),
    .Q(\data_array.data0[3][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12988_ (.CLK(clk),
    .D(_01682_),
    .Q(\data_array.data0[3][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12989_ (.CLK(clk),
    .D(_01683_),
    .Q(\data_array.data0[3][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12990_ (.CLK(clk),
    .D(_01684_),
    .Q(\data_array.data0[3][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12991_ (.CLK(clk),
    .D(_01685_),
    .Q(\data_array.data0[3][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12992_ (.CLK(clk),
    .D(_01686_),
    .Q(\data_array.data0[3][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12993_ (.CLK(clk),
    .D(_01687_),
    .Q(\data_array.data0[3][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12994_ (.CLK(clk),
    .D(_01688_),
    .Q(\data_array.data0[3][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12995_ (.CLK(clk),
    .D(_01689_),
    .Q(\data_array.data0[3][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12996_ (.CLK(clk),
    .D(_01690_),
    .Q(\data_array.data0[3][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12997_ (.CLK(clk),
    .D(_01691_),
    .Q(\data_array.data0[3][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12998_ (.CLK(clk),
    .D(_01692_),
    .Q(\data_array.data0[3][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12999_ (.CLK(clk),
    .D(_01693_),
    .Q(\data_array.data0[3][14] ));
 sky130_fd_sc_hd__dfxtp_2 _13000_ (.CLK(clk),
    .D(_01694_),
    .Q(\data_array.data0[3][15] ));
 sky130_fd_sc_hd__dfxtp_2 _13001_ (.CLK(clk),
    .D(_01695_),
    .Q(\data_array.data0[3][16] ));
 sky130_fd_sc_hd__dfxtp_2 _13002_ (.CLK(clk),
    .D(_01696_),
    .Q(\data_array.data0[3][17] ));
 sky130_fd_sc_hd__dfxtp_2 _13003_ (.CLK(clk),
    .D(_01697_),
    .Q(\data_array.data0[3][18] ));
 sky130_fd_sc_hd__dfxtp_2 _13004_ (.CLK(clk),
    .D(_01698_),
    .Q(\data_array.data0[3][19] ));
 sky130_fd_sc_hd__dfxtp_2 _13005_ (.CLK(clk),
    .D(_01699_),
    .Q(\data_array.data0[3][20] ));
 sky130_fd_sc_hd__dfxtp_2 _13006_ (.CLK(clk),
    .D(_01700_),
    .Q(\data_array.data0[3][21] ));
 sky130_fd_sc_hd__dfxtp_2 _13007_ (.CLK(clk),
    .D(_01701_),
    .Q(\data_array.data0[3][22] ));
 sky130_fd_sc_hd__dfxtp_2 _13008_ (.CLK(clk),
    .D(_01702_),
    .Q(\data_array.data0[3][23] ));
 sky130_fd_sc_hd__dfxtp_2 _13009_ (.CLK(clk),
    .D(_01703_),
    .Q(\data_array.data0[3][24] ));
 sky130_fd_sc_hd__dfxtp_2 _13010_ (.CLK(clk),
    .D(_01704_),
    .Q(\data_array.data0[3][25] ));
 sky130_fd_sc_hd__dfxtp_2 _13011_ (.CLK(clk),
    .D(_01705_),
    .Q(\data_array.data0[3][26] ));
 sky130_fd_sc_hd__dfxtp_2 _13012_ (.CLK(clk),
    .D(_01706_),
    .Q(\data_array.data0[3][27] ));
 sky130_fd_sc_hd__dfxtp_2 _13013_ (.CLK(clk),
    .D(_01707_),
    .Q(\data_array.data0[3][28] ));
 sky130_fd_sc_hd__dfxtp_2 _13014_ (.CLK(clk),
    .D(_01708_),
    .Q(\data_array.data0[3][29] ));
 sky130_fd_sc_hd__dfxtp_2 _13015_ (.CLK(clk),
    .D(_01709_),
    .Q(\data_array.data0[3][30] ));
 sky130_fd_sc_hd__dfxtp_2 _13016_ (.CLK(clk),
    .D(_01710_),
    .Q(\data_array.data0[3][31] ));
 sky130_fd_sc_hd__dfxtp_2 _13017_ (.CLK(clk),
    .D(_01711_),
    .Q(\data_array.data0[3][32] ));
 sky130_fd_sc_hd__dfxtp_2 _13018_ (.CLK(clk),
    .D(_01712_),
    .Q(\data_array.data0[3][33] ));
 sky130_fd_sc_hd__dfxtp_2 _13019_ (.CLK(clk),
    .D(_01713_),
    .Q(\data_array.data0[3][34] ));
 sky130_fd_sc_hd__dfxtp_2 _13020_ (.CLK(clk),
    .D(_01714_),
    .Q(\data_array.data0[3][35] ));
 sky130_fd_sc_hd__dfxtp_2 _13021_ (.CLK(clk),
    .D(_01715_),
    .Q(\data_array.data0[3][36] ));
 sky130_fd_sc_hd__dfxtp_2 _13022_ (.CLK(clk),
    .D(_01716_),
    .Q(\data_array.data0[3][37] ));
 sky130_fd_sc_hd__dfxtp_2 _13023_ (.CLK(clk),
    .D(_01717_),
    .Q(\data_array.data0[3][38] ));
 sky130_fd_sc_hd__dfxtp_2 _13024_ (.CLK(clk),
    .D(_01718_),
    .Q(\data_array.data0[3][39] ));
 sky130_fd_sc_hd__dfxtp_2 _13025_ (.CLK(clk),
    .D(_01719_),
    .Q(\data_array.data0[3][40] ));
 sky130_fd_sc_hd__dfxtp_2 _13026_ (.CLK(clk),
    .D(_01720_),
    .Q(\data_array.data0[3][41] ));
 sky130_fd_sc_hd__dfxtp_2 _13027_ (.CLK(clk),
    .D(_01721_),
    .Q(\data_array.data0[3][42] ));
 sky130_fd_sc_hd__dfxtp_2 _13028_ (.CLK(clk),
    .D(_01722_),
    .Q(\data_array.data0[3][43] ));
 sky130_fd_sc_hd__dfxtp_2 _13029_ (.CLK(clk),
    .D(_01723_),
    .Q(\data_array.data0[3][44] ));
 sky130_fd_sc_hd__dfxtp_2 _13030_ (.CLK(clk),
    .D(_01724_),
    .Q(\data_array.data0[3][45] ));
 sky130_fd_sc_hd__dfxtp_2 _13031_ (.CLK(clk),
    .D(_01725_),
    .Q(\data_array.data0[3][46] ));
 sky130_fd_sc_hd__dfxtp_2 _13032_ (.CLK(clk),
    .D(_01726_),
    .Q(\data_array.data0[3][47] ));
 sky130_fd_sc_hd__dfxtp_2 _13033_ (.CLK(clk),
    .D(_01727_),
    .Q(\data_array.data0[3][48] ));
 sky130_fd_sc_hd__dfxtp_2 _13034_ (.CLK(clk),
    .D(_01728_),
    .Q(\data_array.data0[3][49] ));
 sky130_fd_sc_hd__dfxtp_2 _13035_ (.CLK(clk),
    .D(_01729_),
    .Q(\data_array.data0[3][50] ));
 sky130_fd_sc_hd__dfxtp_2 _13036_ (.CLK(clk),
    .D(_01730_),
    .Q(\data_array.data0[3][51] ));
 sky130_fd_sc_hd__dfxtp_2 _13037_ (.CLK(clk),
    .D(_01731_),
    .Q(\data_array.data0[3][52] ));
 sky130_fd_sc_hd__dfxtp_2 _13038_ (.CLK(clk),
    .D(_01732_),
    .Q(\data_array.data0[3][53] ));
 sky130_fd_sc_hd__dfxtp_2 _13039_ (.CLK(clk),
    .D(_01733_),
    .Q(\data_array.data0[3][54] ));
 sky130_fd_sc_hd__dfxtp_2 _13040_ (.CLK(clk),
    .D(_01734_),
    .Q(\data_array.data0[3][55] ));
 sky130_fd_sc_hd__dfxtp_2 _13041_ (.CLK(clk),
    .D(_01735_),
    .Q(\data_array.data0[3][56] ));
 sky130_fd_sc_hd__dfxtp_2 _13042_ (.CLK(clk),
    .D(_01736_),
    .Q(\data_array.data0[3][57] ));
 sky130_fd_sc_hd__dfxtp_2 _13043_ (.CLK(clk),
    .D(_01737_),
    .Q(\data_array.data0[3][58] ));
 sky130_fd_sc_hd__dfxtp_2 _13044_ (.CLK(clk),
    .D(_01738_),
    .Q(\data_array.data0[3][59] ));
 sky130_fd_sc_hd__dfxtp_2 _13045_ (.CLK(clk),
    .D(_01739_),
    .Q(\data_array.data0[3][60] ));
 sky130_fd_sc_hd__dfxtp_2 _13046_ (.CLK(clk),
    .D(_01740_),
    .Q(\data_array.data0[3][61] ));
 sky130_fd_sc_hd__dfxtp_2 _13047_ (.CLK(clk),
    .D(_01741_),
    .Q(\data_array.data0[3][62] ));
 sky130_fd_sc_hd__dfxtp_2 _13048_ (.CLK(clk),
    .D(_01742_),
    .Q(\data_array.data0[3][63] ));
 sky130_fd_sc_hd__dfxtp_2 _13049_ (.CLK(clk),
    .D(_01743_),
    .Q(\data_array.data1[13][0] ));
 sky130_fd_sc_hd__dfxtp_2 _13050_ (.CLK(clk),
    .D(_01744_),
    .Q(\data_array.data1[13][1] ));
 sky130_fd_sc_hd__dfxtp_2 _13051_ (.CLK(clk),
    .D(_01745_),
    .Q(\data_array.data1[13][2] ));
 sky130_fd_sc_hd__dfxtp_2 _13052_ (.CLK(clk),
    .D(_01746_),
    .Q(\data_array.data1[13][3] ));
 sky130_fd_sc_hd__dfxtp_2 _13053_ (.CLK(clk),
    .D(_01747_),
    .Q(\data_array.data1[13][4] ));
 sky130_fd_sc_hd__dfxtp_2 _13054_ (.CLK(clk),
    .D(_01748_),
    .Q(\data_array.data1[13][5] ));
 sky130_fd_sc_hd__dfxtp_2 _13055_ (.CLK(clk),
    .D(_01749_),
    .Q(\data_array.data1[13][6] ));
 sky130_fd_sc_hd__dfxtp_2 _13056_ (.CLK(clk),
    .D(_01750_),
    .Q(\data_array.data1[13][7] ));
 sky130_fd_sc_hd__dfxtp_2 _13057_ (.CLK(clk),
    .D(_01751_),
    .Q(\data_array.data1[13][8] ));
 sky130_fd_sc_hd__dfxtp_2 _13058_ (.CLK(clk),
    .D(_01752_),
    .Q(\data_array.data1[13][9] ));
 sky130_fd_sc_hd__dfxtp_2 _13059_ (.CLK(clk),
    .D(_01753_),
    .Q(\data_array.data1[13][10] ));
 sky130_fd_sc_hd__dfxtp_2 _13060_ (.CLK(clk),
    .D(_01754_),
    .Q(\data_array.data1[13][11] ));
 sky130_fd_sc_hd__dfxtp_2 _13061_ (.CLK(clk),
    .D(_01755_),
    .Q(\data_array.data1[13][12] ));
 sky130_fd_sc_hd__dfxtp_2 _13062_ (.CLK(clk),
    .D(_01756_),
    .Q(\data_array.data1[13][13] ));
 sky130_fd_sc_hd__dfxtp_2 _13063_ (.CLK(clk),
    .D(_01757_),
    .Q(\data_array.data1[13][14] ));
 sky130_fd_sc_hd__dfxtp_2 _13064_ (.CLK(clk),
    .D(_01758_),
    .Q(\data_array.data1[13][15] ));
 sky130_fd_sc_hd__dfxtp_2 _13065_ (.CLK(clk),
    .D(_01759_),
    .Q(\data_array.data1[13][16] ));
 sky130_fd_sc_hd__dfxtp_2 _13066_ (.CLK(clk),
    .D(_01760_),
    .Q(\data_array.data1[13][17] ));
 sky130_fd_sc_hd__dfxtp_2 _13067_ (.CLK(clk),
    .D(_01761_),
    .Q(\data_array.data1[13][18] ));
 sky130_fd_sc_hd__dfxtp_2 _13068_ (.CLK(clk),
    .D(_01762_),
    .Q(\data_array.data1[13][19] ));
 sky130_fd_sc_hd__dfxtp_2 _13069_ (.CLK(clk),
    .D(_01763_),
    .Q(\data_array.data1[13][20] ));
 sky130_fd_sc_hd__dfxtp_2 _13070_ (.CLK(clk),
    .D(_01764_),
    .Q(\data_array.data1[13][21] ));
 sky130_fd_sc_hd__dfxtp_2 _13071_ (.CLK(clk),
    .D(_01765_),
    .Q(\data_array.data1[13][22] ));
 sky130_fd_sc_hd__dfxtp_2 _13072_ (.CLK(clk),
    .D(_01766_),
    .Q(\data_array.data1[13][23] ));
 sky130_fd_sc_hd__dfxtp_2 _13073_ (.CLK(clk),
    .D(_01767_),
    .Q(\data_array.data1[13][24] ));
 sky130_fd_sc_hd__dfxtp_2 _13074_ (.CLK(clk),
    .D(_01768_),
    .Q(\data_array.data1[13][25] ));
 sky130_fd_sc_hd__dfxtp_2 _13075_ (.CLK(clk),
    .D(_01769_),
    .Q(\data_array.data1[13][26] ));
 sky130_fd_sc_hd__dfxtp_2 _13076_ (.CLK(clk),
    .D(_01770_),
    .Q(\data_array.data1[13][27] ));
 sky130_fd_sc_hd__dfxtp_2 _13077_ (.CLK(clk),
    .D(_01771_),
    .Q(\data_array.data1[13][28] ));
 sky130_fd_sc_hd__dfxtp_2 _13078_ (.CLK(clk),
    .D(_01772_),
    .Q(\data_array.data1[13][29] ));
 sky130_fd_sc_hd__dfxtp_2 _13079_ (.CLK(clk),
    .D(_01773_),
    .Q(\data_array.data1[13][30] ));
 sky130_fd_sc_hd__dfxtp_2 _13080_ (.CLK(clk),
    .D(_01774_),
    .Q(\data_array.data1[13][31] ));
 sky130_fd_sc_hd__dfxtp_2 _13081_ (.CLK(clk),
    .D(_01775_),
    .Q(\data_array.data1[13][32] ));
 sky130_fd_sc_hd__dfxtp_2 _13082_ (.CLK(clk),
    .D(_01776_),
    .Q(\data_array.data1[13][33] ));
 sky130_fd_sc_hd__dfxtp_2 _13083_ (.CLK(clk),
    .D(_01777_),
    .Q(\data_array.data1[13][34] ));
 sky130_fd_sc_hd__dfxtp_2 _13084_ (.CLK(clk),
    .D(_01778_),
    .Q(\data_array.data1[13][35] ));
 sky130_fd_sc_hd__dfxtp_2 _13085_ (.CLK(clk),
    .D(_01779_),
    .Q(\data_array.data1[13][36] ));
 sky130_fd_sc_hd__dfxtp_2 _13086_ (.CLK(clk),
    .D(_01780_),
    .Q(\data_array.data1[13][37] ));
 sky130_fd_sc_hd__dfxtp_2 _13087_ (.CLK(clk),
    .D(_01781_),
    .Q(\data_array.data1[13][38] ));
 sky130_fd_sc_hd__dfxtp_2 _13088_ (.CLK(clk),
    .D(_01782_),
    .Q(\data_array.data1[13][39] ));
 sky130_fd_sc_hd__dfxtp_2 _13089_ (.CLK(clk),
    .D(_01783_),
    .Q(\data_array.data1[13][40] ));
 sky130_fd_sc_hd__dfxtp_2 _13090_ (.CLK(clk),
    .D(_01784_),
    .Q(\data_array.data1[13][41] ));
 sky130_fd_sc_hd__dfxtp_2 _13091_ (.CLK(clk),
    .D(_01785_),
    .Q(\data_array.data1[13][42] ));
 sky130_fd_sc_hd__dfxtp_2 _13092_ (.CLK(clk),
    .D(_01786_),
    .Q(\data_array.data1[13][43] ));
 sky130_fd_sc_hd__dfxtp_2 _13093_ (.CLK(clk),
    .D(_01787_),
    .Q(\data_array.data1[13][44] ));
 sky130_fd_sc_hd__dfxtp_2 _13094_ (.CLK(clk),
    .D(_01788_),
    .Q(\data_array.data1[13][45] ));
 sky130_fd_sc_hd__dfxtp_2 _13095_ (.CLK(clk),
    .D(_01789_),
    .Q(\data_array.data1[13][46] ));
 sky130_fd_sc_hd__dfxtp_2 _13096_ (.CLK(clk),
    .D(_01790_),
    .Q(\data_array.data1[13][47] ));
 sky130_fd_sc_hd__dfxtp_2 _13097_ (.CLK(clk),
    .D(_01791_),
    .Q(\data_array.data1[13][48] ));
 sky130_fd_sc_hd__dfxtp_2 _13098_ (.CLK(clk),
    .D(_01792_),
    .Q(\data_array.data1[13][49] ));
 sky130_fd_sc_hd__dfxtp_2 _13099_ (.CLK(clk),
    .D(_01793_),
    .Q(\data_array.data1[13][50] ));
 sky130_fd_sc_hd__dfxtp_2 _13100_ (.CLK(clk),
    .D(_01794_),
    .Q(\data_array.data1[13][51] ));
 sky130_fd_sc_hd__dfxtp_2 _13101_ (.CLK(clk),
    .D(_01795_),
    .Q(\data_array.data1[13][52] ));
 sky130_fd_sc_hd__dfxtp_2 _13102_ (.CLK(clk),
    .D(_01796_),
    .Q(\data_array.data1[13][53] ));
 sky130_fd_sc_hd__dfxtp_2 _13103_ (.CLK(clk),
    .D(_01797_),
    .Q(\data_array.data1[13][54] ));
 sky130_fd_sc_hd__dfxtp_2 _13104_ (.CLK(clk),
    .D(_01798_),
    .Q(\data_array.data1[13][55] ));
 sky130_fd_sc_hd__dfxtp_2 _13105_ (.CLK(clk),
    .D(_01799_),
    .Q(\data_array.data1[13][56] ));
 sky130_fd_sc_hd__dfxtp_2 _13106_ (.CLK(clk),
    .D(_01800_),
    .Q(\data_array.data1[13][57] ));
 sky130_fd_sc_hd__dfxtp_2 _13107_ (.CLK(clk),
    .D(_01801_),
    .Q(\data_array.data1[13][58] ));
 sky130_fd_sc_hd__dfxtp_2 _13108_ (.CLK(clk),
    .D(_01802_),
    .Q(\data_array.data1[13][59] ));
 sky130_fd_sc_hd__dfxtp_2 _13109_ (.CLK(clk),
    .D(_01803_),
    .Q(\data_array.data1[13][60] ));
 sky130_fd_sc_hd__dfxtp_2 _13110_ (.CLK(clk),
    .D(_01804_),
    .Q(\data_array.data1[13][61] ));
 sky130_fd_sc_hd__dfxtp_2 _13111_ (.CLK(clk),
    .D(_01805_),
    .Q(\data_array.data1[13][62] ));
 sky130_fd_sc_hd__dfxtp_2 _13112_ (.CLK(clk),
    .D(_01806_),
    .Q(\data_array.data1[13][63] ));
 sky130_fd_sc_hd__dfxtp_2 _13113_ (.CLK(clk),
    .D(_01807_),
    .Q(\tag_array.tag0[3][0] ));
 sky130_fd_sc_hd__dfxtp_2 _13114_ (.CLK(clk),
    .D(_01808_),
    .Q(\tag_array.tag0[3][1] ));
 sky130_fd_sc_hd__dfxtp_2 _13115_ (.CLK(clk),
    .D(_01809_),
    .Q(\tag_array.tag0[3][2] ));
 sky130_fd_sc_hd__dfxtp_2 _13116_ (.CLK(clk),
    .D(_01810_),
    .Q(\tag_array.tag0[3][3] ));
 sky130_fd_sc_hd__dfxtp_2 _13117_ (.CLK(clk),
    .D(_01811_),
    .Q(\tag_array.tag0[3][4] ));
 sky130_fd_sc_hd__dfxtp_2 _13118_ (.CLK(clk),
    .D(_01812_),
    .Q(\tag_array.tag0[3][5] ));
 sky130_fd_sc_hd__dfxtp_2 _13119_ (.CLK(clk),
    .D(_01813_),
    .Q(\tag_array.tag0[3][6] ));
 sky130_fd_sc_hd__dfxtp_2 _13120_ (.CLK(clk),
    .D(_01814_),
    .Q(\tag_array.tag0[3][7] ));
 sky130_fd_sc_hd__dfxtp_2 _13121_ (.CLK(clk),
    .D(_01815_),
    .Q(\tag_array.tag0[3][8] ));
 sky130_fd_sc_hd__dfxtp_2 _13122_ (.CLK(clk),
    .D(_01816_),
    .Q(\tag_array.tag0[3][9] ));
 sky130_fd_sc_hd__dfxtp_2 _13123_ (.CLK(clk),
    .D(_01817_),
    .Q(\tag_array.tag0[3][10] ));
 sky130_fd_sc_hd__dfxtp_2 _13124_ (.CLK(clk),
    .D(_01818_),
    .Q(\tag_array.tag0[3][11] ));
 sky130_fd_sc_hd__dfxtp_2 _13125_ (.CLK(clk),
    .D(_01819_),
    .Q(\tag_array.tag0[3][12] ));
 sky130_fd_sc_hd__dfxtp_2 _13126_ (.CLK(clk),
    .D(_01820_),
    .Q(\tag_array.tag0[3][13] ));
 sky130_fd_sc_hd__dfxtp_2 _13127_ (.CLK(clk),
    .D(_01821_),
    .Q(\tag_array.tag0[3][14] ));
 sky130_fd_sc_hd__dfxtp_2 _13128_ (.CLK(clk),
    .D(_01822_),
    .Q(\tag_array.tag0[3][15] ));
 sky130_fd_sc_hd__dfxtp_2 _13129_ (.CLK(clk),
    .D(_01823_),
    .Q(\tag_array.tag0[3][16] ));
 sky130_fd_sc_hd__dfxtp_2 _13130_ (.CLK(clk),
    .D(_01824_),
    .Q(\tag_array.tag0[3][17] ));
 sky130_fd_sc_hd__dfxtp_2 _13131_ (.CLK(clk),
    .D(_01825_),
    .Q(\tag_array.tag0[3][18] ));
 sky130_fd_sc_hd__dfxtp_2 _13132_ (.CLK(clk),
    .D(_01826_),
    .Q(\tag_array.tag0[3][19] ));
 sky130_fd_sc_hd__dfxtp_2 _13133_ (.CLK(clk),
    .D(_01827_),
    .Q(\tag_array.tag0[3][20] ));
 sky130_fd_sc_hd__dfxtp_2 _13134_ (.CLK(clk),
    .D(_01828_),
    .Q(\tag_array.tag0[3][21] ));
 sky130_fd_sc_hd__dfxtp_2 _13135_ (.CLK(clk),
    .D(_01829_),
    .Q(\tag_array.tag0[3][22] ));
 sky130_fd_sc_hd__dfxtp_2 _13136_ (.CLK(clk),
    .D(_01830_),
    .Q(\tag_array.tag0[3][23] ));
 sky130_fd_sc_hd__dfxtp_2 _13137_ (.CLK(clk),
    .D(_01831_),
    .Q(\tag_array.tag0[3][24] ));
 sky130_fd_sc_hd__dfxtp_2 _13138_ (.CLK(clk),
    .D(_01832_),
    .Q(\tag_array.tag1[8][0] ));
 sky130_fd_sc_hd__dfxtp_2 _13139_ (.CLK(clk),
    .D(_01833_),
    .Q(\tag_array.tag1[8][1] ));
 sky130_fd_sc_hd__dfxtp_2 _13140_ (.CLK(clk),
    .D(_01834_),
    .Q(\tag_array.tag1[8][2] ));
 sky130_fd_sc_hd__dfxtp_2 _13141_ (.CLK(clk),
    .D(_01835_),
    .Q(\tag_array.tag1[8][3] ));
 sky130_fd_sc_hd__dfxtp_2 _13142_ (.CLK(clk),
    .D(_01836_),
    .Q(\tag_array.tag1[8][4] ));
 sky130_fd_sc_hd__dfxtp_2 _13143_ (.CLK(clk),
    .D(_01837_),
    .Q(\tag_array.tag1[8][5] ));
 sky130_fd_sc_hd__dfxtp_2 _13144_ (.CLK(clk),
    .D(_01838_),
    .Q(\tag_array.tag1[8][6] ));
 sky130_fd_sc_hd__dfxtp_2 _13145_ (.CLK(clk),
    .D(_01839_),
    .Q(\tag_array.tag1[8][7] ));
 sky130_fd_sc_hd__dfxtp_2 _13146_ (.CLK(clk),
    .D(_01840_),
    .Q(\tag_array.tag1[8][8] ));
 sky130_fd_sc_hd__dfxtp_2 _13147_ (.CLK(clk),
    .D(_01841_),
    .Q(\tag_array.tag1[8][9] ));
 sky130_fd_sc_hd__dfxtp_2 _13148_ (.CLK(clk),
    .D(_01842_),
    .Q(\tag_array.tag1[8][10] ));
 sky130_fd_sc_hd__dfxtp_2 _13149_ (.CLK(clk),
    .D(_01843_),
    .Q(\tag_array.tag1[8][11] ));
 sky130_fd_sc_hd__dfxtp_2 _13150_ (.CLK(clk),
    .D(_01844_),
    .Q(\tag_array.tag1[8][12] ));
 sky130_fd_sc_hd__dfxtp_2 _13151_ (.CLK(clk),
    .D(_01845_),
    .Q(\tag_array.tag1[8][13] ));
 sky130_fd_sc_hd__dfxtp_2 _13152_ (.CLK(clk),
    .D(_01846_),
    .Q(\tag_array.tag1[8][14] ));
 sky130_fd_sc_hd__dfxtp_2 _13153_ (.CLK(clk),
    .D(_01847_),
    .Q(\tag_array.tag1[8][15] ));
 sky130_fd_sc_hd__dfxtp_2 _13154_ (.CLK(clk),
    .D(_01848_),
    .Q(\tag_array.tag1[8][16] ));
 sky130_fd_sc_hd__dfxtp_2 _13155_ (.CLK(clk),
    .D(_01849_),
    .Q(\tag_array.tag1[8][17] ));
 sky130_fd_sc_hd__dfxtp_2 _13156_ (.CLK(clk),
    .D(_01850_),
    .Q(\tag_array.tag1[8][18] ));
 sky130_fd_sc_hd__dfxtp_2 _13157_ (.CLK(clk),
    .D(_01851_),
    .Q(\tag_array.tag1[8][19] ));
 sky130_fd_sc_hd__dfxtp_2 _13158_ (.CLK(clk),
    .D(_01852_),
    .Q(\tag_array.tag1[8][20] ));
 sky130_fd_sc_hd__dfxtp_2 _13159_ (.CLK(clk),
    .D(_01853_),
    .Q(\tag_array.tag1[8][21] ));
 sky130_fd_sc_hd__dfxtp_2 _13160_ (.CLK(clk),
    .D(_01854_),
    .Q(\tag_array.tag1[8][22] ));
 sky130_fd_sc_hd__dfxtp_2 _13161_ (.CLK(clk),
    .D(_01855_),
    .Q(\tag_array.tag1[8][23] ));
 sky130_fd_sc_hd__dfxtp_2 _13162_ (.CLK(clk),
    .D(_01856_),
    .Q(\tag_array.tag1[8][24] ));
 sky130_fd_sc_hd__dfxtp_2 _13163_ (.CLK(clk),
    .D(_00064_),
    .Q(\data_array.rdata1[0] ));
 sky130_fd_sc_hd__dfxtp_2 _13164_ (.CLK(clk),
    .D(_00075_),
    .Q(\data_array.rdata1[1] ));
 sky130_fd_sc_hd__dfxtp_2 _13165_ (.CLK(clk),
    .D(_00086_),
    .Q(\data_array.rdata1[2] ));
 sky130_fd_sc_hd__dfxtp_2 _13166_ (.CLK(clk),
    .D(_00097_),
    .Q(\data_array.rdata1[3] ));
 sky130_fd_sc_hd__dfxtp_2 _13167_ (.CLK(clk),
    .D(_00108_),
    .Q(\data_array.rdata1[4] ));
 sky130_fd_sc_hd__dfxtp_2 _13168_ (.CLK(clk),
    .D(_00119_),
    .Q(\data_array.rdata1[5] ));
 sky130_fd_sc_hd__dfxtp_2 _13169_ (.CLK(clk),
    .D(_00124_),
    .Q(\data_array.rdata1[6] ));
 sky130_fd_sc_hd__dfxtp_2 _13170_ (.CLK(clk),
    .D(_00125_),
    .Q(\data_array.rdata1[7] ));
 sky130_fd_sc_hd__dfxtp_2 _13171_ (.CLK(clk),
    .D(_00126_),
    .Q(\data_array.rdata1[8] ));
 sky130_fd_sc_hd__dfxtp_2 _13172_ (.CLK(clk),
    .D(_00127_),
    .Q(\data_array.rdata1[9] ));
 sky130_fd_sc_hd__dfxtp_2 _13173_ (.CLK(clk),
    .D(_00065_),
    .Q(\data_array.rdata1[10] ));
 sky130_fd_sc_hd__dfxtp_2 _13174_ (.CLK(clk),
    .D(_00066_),
    .Q(\data_array.rdata1[11] ));
 sky130_fd_sc_hd__dfxtp_2 _13175_ (.CLK(clk),
    .D(_00067_),
    .Q(\data_array.rdata1[12] ));
 sky130_fd_sc_hd__dfxtp_2 _13176_ (.CLK(clk),
    .D(_00068_),
    .Q(\data_array.rdata1[13] ));
 sky130_fd_sc_hd__dfxtp_2 _13177_ (.CLK(clk),
    .D(_00069_),
    .Q(\data_array.rdata1[14] ));
 sky130_fd_sc_hd__dfxtp_2 _13178_ (.CLK(clk),
    .D(_00070_),
    .Q(\data_array.rdata1[15] ));
 sky130_fd_sc_hd__dfxtp_2 _13179_ (.CLK(clk),
    .D(_00071_),
    .Q(\data_array.rdata1[16] ));
 sky130_fd_sc_hd__dfxtp_2 _13180_ (.CLK(clk),
    .D(_00072_),
    .Q(\data_array.rdata1[17] ));
 sky130_fd_sc_hd__dfxtp_2 _13181_ (.CLK(clk),
    .D(_00073_),
    .Q(\data_array.rdata1[18] ));
 sky130_fd_sc_hd__dfxtp_2 _13182_ (.CLK(clk),
    .D(_00074_),
    .Q(\data_array.rdata1[19] ));
 sky130_fd_sc_hd__dfxtp_2 _13183_ (.CLK(clk),
    .D(_00076_),
    .Q(\data_array.rdata1[20] ));
 sky130_fd_sc_hd__dfxtp_2 _13184_ (.CLK(clk),
    .D(_00077_),
    .Q(\data_array.rdata1[21] ));
 sky130_fd_sc_hd__dfxtp_2 _13185_ (.CLK(clk),
    .D(_00078_),
    .Q(\data_array.rdata1[22] ));
 sky130_fd_sc_hd__dfxtp_2 _13186_ (.CLK(clk),
    .D(_00079_),
    .Q(\data_array.rdata1[23] ));
 sky130_fd_sc_hd__dfxtp_2 _13187_ (.CLK(clk),
    .D(_00080_),
    .Q(\data_array.rdata1[24] ));
 sky130_fd_sc_hd__dfxtp_2 _13188_ (.CLK(clk),
    .D(_00081_),
    .Q(\data_array.rdata1[25] ));
 sky130_fd_sc_hd__dfxtp_2 _13189_ (.CLK(clk),
    .D(_00082_),
    .Q(\data_array.rdata1[26] ));
 sky130_fd_sc_hd__dfxtp_2 _13190_ (.CLK(clk),
    .D(_00083_),
    .Q(\data_array.rdata1[27] ));
 sky130_fd_sc_hd__dfxtp_2 _13191_ (.CLK(clk),
    .D(_00084_),
    .Q(\data_array.rdata1[28] ));
 sky130_fd_sc_hd__dfxtp_2 _13192_ (.CLK(clk),
    .D(_00085_),
    .Q(\data_array.rdata1[29] ));
 sky130_fd_sc_hd__dfxtp_2 _13193_ (.CLK(clk),
    .D(_00087_),
    .Q(\data_array.rdata1[30] ));
 sky130_fd_sc_hd__dfxtp_2 _13194_ (.CLK(clk),
    .D(_00088_),
    .Q(\data_array.rdata1[31] ));
 sky130_fd_sc_hd__dfxtp_2 _13195_ (.CLK(clk),
    .D(_00089_),
    .Q(\data_array.rdata1[32] ));
 sky130_fd_sc_hd__dfxtp_2 _13196_ (.CLK(clk),
    .D(_00090_),
    .Q(\data_array.rdata1[33] ));
 sky130_fd_sc_hd__dfxtp_2 _13197_ (.CLK(clk),
    .D(_00091_),
    .Q(\data_array.rdata1[34] ));
 sky130_fd_sc_hd__dfxtp_2 _13198_ (.CLK(clk),
    .D(_00092_),
    .Q(\data_array.rdata1[35] ));
 sky130_fd_sc_hd__dfxtp_2 _13199_ (.CLK(clk),
    .D(_00093_),
    .Q(\data_array.rdata1[36] ));
 sky130_fd_sc_hd__dfxtp_2 _13200_ (.CLK(clk),
    .D(_00094_),
    .Q(\data_array.rdata1[37] ));
 sky130_fd_sc_hd__dfxtp_2 _13201_ (.CLK(clk),
    .D(_00095_),
    .Q(\data_array.rdata1[38] ));
 sky130_fd_sc_hd__dfxtp_2 _13202_ (.CLK(clk),
    .D(_00096_),
    .Q(\data_array.rdata1[39] ));
 sky130_fd_sc_hd__dfxtp_2 _13203_ (.CLK(clk),
    .D(_00098_),
    .Q(\data_array.rdata1[40] ));
 sky130_fd_sc_hd__dfxtp_2 _13204_ (.CLK(clk),
    .D(_00099_),
    .Q(\data_array.rdata1[41] ));
 sky130_fd_sc_hd__dfxtp_2 _13205_ (.CLK(clk),
    .D(_00100_),
    .Q(\data_array.rdata1[42] ));
 sky130_fd_sc_hd__dfxtp_2 _13206_ (.CLK(clk),
    .D(_00101_),
    .Q(\data_array.rdata1[43] ));
 sky130_fd_sc_hd__dfxtp_2 _13207_ (.CLK(clk),
    .D(_00102_),
    .Q(\data_array.rdata1[44] ));
 sky130_fd_sc_hd__dfxtp_2 _13208_ (.CLK(clk),
    .D(_00103_),
    .Q(\data_array.rdata1[45] ));
 sky130_fd_sc_hd__dfxtp_2 _13209_ (.CLK(clk),
    .D(_00104_),
    .Q(\data_array.rdata1[46] ));
 sky130_fd_sc_hd__dfxtp_2 _13210_ (.CLK(clk),
    .D(_00105_),
    .Q(\data_array.rdata1[47] ));
 sky130_fd_sc_hd__dfxtp_2 _13211_ (.CLK(clk),
    .D(_00106_),
    .Q(\data_array.rdata1[48] ));
 sky130_fd_sc_hd__dfxtp_2 _13212_ (.CLK(clk),
    .D(_00107_),
    .Q(\data_array.rdata1[49] ));
 sky130_fd_sc_hd__dfxtp_2 _13213_ (.CLK(clk),
    .D(_00109_),
    .Q(\data_array.rdata1[50] ));
 sky130_fd_sc_hd__dfxtp_2 _13214_ (.CLK(clk),
    .D(_00110_),
    .Q(\data_array.rdata1[51] ));
 sky130_fd_sc_hd__dfxtp_2 _13215_ (.CLK(clk),
    .D(_00111_),
    .Q(\data_array.rdata1[52] ));
 sky130_fd_sc_hd__dfxtp_2 _13216_ (.CLK(clk),
    .D(_00112_),
    .Q(\data_array.rdata1[53] ));
 sky130_fd_sc_hd__dfxtp_2 _13217_ (.CLK(clk),
    .D(_00113_),
    .Q(\data_array.rdata1[54] ));
 sky130_fd_sc_hd__dfxtp_2 _13218_ (.CLK(clk),
    .D(_00114_),
    .Q(\data_array.rdata1[55] ));
 sky130_fd_sc_hd__dfxtp_2 _13219_ (.CLK(clk),
    .D(_00115_),
    .Q(\data_array.rdata1[56] ));
 sky130_fd_sc_hd__dfxtp_2 _13220_ (.CLK(clk),
    .D(_00116_),
    .Q(\data_array.rdata1[57] ));
 sky130_fd_sc_hd__dfxtp_2 _13221_ (.CLK(clk),
    .D(_00117_),
    .Q(\data_array.rdata1[58] ));
 sky130_fd_sc_hd__dfxtp_2 _13222_ (.CLK(clk),
    .D(_00118_),
    .Q(\data_array.rdata1[59] ));
 sky130_fd_sc_hd__dfxtp_2 _13223_ (.CLK(clk),
    .D(_00120_),
    .Q(\data_array.rdata1[60] ));
 sky130_fd_sc_hd__dfxtp_2 _13224_ (.CLK(clk),
    .D(_00121_),
    .Q(\data_array.rdata1[61] ));
 sky130_fd_sc_hd__dfxtp_2 _13225_ (.CLK(clk),
    .D(_00122_),
    .Q(\data_array.rdata1[62] ));
 sky130_fd_sc_hd__dfxtp_2 _13226_ (.CLK(clk),
    .D(_00123_),
    .Q(\data_array.rdata1[63] ));
 sky130_fd_sc_hd__dfxtp_2 _13227_ (.CLK(clk),
    .D(_01857_),
    .Q(\data_array.data0[11][0] ));
 sky130_fd_sc_hd__dfxtp_2 _13228_ (.CLK(clk),
    .D(_01858_),
    .Q(\data_array.data0[11][1] ));
 sky130_fd_sc_hd__dfxtp_2 _13229_ (.CLK(clk),
    .D(_01859_),
    .Q(\data_array.data0[11][2] ));
 sky130_fd_sc_hd__dfxtp_2 _13230_ (.CLK(clk),
    .D(_01860_),
    .Q(\data_array.data0[11][3] ));
 sky130_fd_sc_hd__dfxtp_2 _13231_ (.CLK(clk),
    .D(_01861_),
    .Q(\data_array.data0[11][4] ));
 sky130_fd_sc_hd__dfxtp_2 _13232_ (.CLK(clk),
    .D(_01862_),
    .Q(\data_array.data0[11][5] ));
 sky130_fd_sc_hd__dfxtp_2 _13233_ (.CLK(clk),
    .D(_01863_),
    .Q(\data_array.data0[11][6] ));
 sky130_fd_sc_hd__dfxtp_2 _13234_ (.CLK(clk),
    .D(_01864_),
    .Q(\data_array.data0[11][7] ));
 sky130_fd_sc_hd__dfxtp_2 _13235_ (.CLK(clk),
    .D(_01865_),
    .Q(\data_array.data0[11][8] ));
 sky130_fd_sc_hd__dfxtp_2 _13236_ (.CLK(clk),
    .D(_01866_),
    .Q(\data_array.data0[11][9] ));
 sky130_fd_sc_hd__dfxtp_2 _13237_ (.CLK(clk),
    .D(_01867_),
    .Q(\data_array.data0[11][10] ));
 sky130_fd_sc_hd__dfxtp_2 _13238_ (.CLK(clk),
    .D(_01868_),
    .Q(\data_array.data0[11][11] ));
 sky130_fd_sc_hd__dfxtp_2 _13239_ (.CLK(clk),
    .D(_01869_),
    .Q(\data_array.data0[11][12] ));
 sky130_fd_sc_hd__dfxtp_2 _13240_ (.CLK(clk),
    .D(_01870_),
    .Q(\data_array.data0[11][13] ));
 sky130_fd_sc_hd__dfxtp_2 _13241_ (.CLK(clk),
    .D(_01871_),
    .Q(\data_array.data0[11][14] ));
 sky130_fd_sc_hd__dfxtp_2 _13242_ (.CLK(clk),
    .D(_01872_),
    .Q(\data_array.data0[11][15] ));
 sky130_fd_sc_hd__dfxtp_2 _13243_ (.CLK(clk),
    .D(_01873_),
    .Q(\data_array.data0[11][16] ));
 sky130_fd_sc_hd__dfxtp_2 _13244_ (.CLK(clk),
    .D(_01874_),
    .Q(\data_array.data0[11][17] ));
 sky130_fd_sc_hd__dfxtp_2 _13245_ (.CLK(clk),
    .D(_01875_),
    .Q(\data_array.data0[11][18] ));
 sky130_fd_sc_hd__dfxtp_2 _13246_ (.CLK(clk),
    .D(_01876_),
    .Q(\data_array.data0[11][19] ));
 sky130_fd_sc_hd__dfxtp_2 _13247_ (.CLK(clk),
    .D(_01877_),
    .Q(\data_array.data0[11][20] ));
 sky130_fd_sc_hd__dfxtp_2 _13248_ (.CLK(clk),
    .D(_01878_),
    .Q(\data_array.data0[11][21] ));
 sky130_fd_sc_hd__dfxtp_2 _13249_ (.CLK(clk),
    .D(_01879_),
    .Q(\data_array.data0[11][22] ));
 sky130_fd_sc_hd__dfxtp_2 _13250_ (.CLK(clk),
    .D(_01880_),
    .Q(\data_array.data0[11][23] ));
 sky130_fd_sc_hd__dfxtp_2 _13251_ (.CLK(clk),
    .D(_01881_),
    .Q(\data_array.data0[11][24] ));
 sky130_fd_sc_hd__dfxtp_2 _13252_ (.CLK(clk),
    .D(_01882_),
    .Q(\data_array.data0[11][25] ));
 sky130_fd_sc_hd__dfxtp_2 _13253_ (.CLK(clk),
    .D(_01883_),
    .Q(\data_array.data0[11][26] ));
 sky130_fd_sc_hd__dfxtp_2 _13254_ (.CLK(clk),
    .D(_01884_),
    .Q(\data_array.data0[11][27] ));
 sky130_fd_sc_hd__dfxtp_2 _13255_ (.CLK(clk),
    .D(_01885_),
    .Q(\data_array.data0[11][28] ));
 sky130_fd_sc_hd__dfxtp_2 _13256_ (.CLK(clk),
    .D(_01886_),
    .Q(\data_array.data0[11][29] ));
 sky130_fd_sc_hd__dfxtp_2 _13257_ (.CLK(clk),
    .D(_01887_),
    .Q(\data_array.data0[11][30] ));
 sky130_fd_sc_hd__dfxtp_2 _13258_ (.CLK(clk),
    .D(_01888_),
    .Q(\data_array.data0[11][31] ));
 sky130_fd_sc_hd__dfxtp_2 _13259_ (.CLK(clk),
    .D(_01889_),
    .Q(\data_array.data0[11][32] ));
 sky130_fd_sc_hd__dfxtp_2 _13260_ (.CLK(clk),
    .D(_01890_),
    .Q(\data_array.data0[11][33] ));
 sky130_fd_sc_hd__dfxtp_2 _13261_ (.CLK(clk),
    .D(_01891_),
    .Q(\data_array.data0[11][34] ));
 sky130_fd_sc_hd__dfxtp_2 _13262_ (.CLK(clk),
    .D(_01892_),
    .Q(\data_array.data0[11][35] ));
 sky130_fd_sc_hd__dfxtp_2 _13263_ (.CLK(clk),
    .D(_01893_),
    .Q(\data_array.data0[11][36] ));
 sky130_fd_sc_hd__dfxtp_2 _13264_ (.CLK(clk),
    .D(_01894_),
    .Q(\data_array.data0[11][37] ));
 sky130_fd_sc_hd__dfxtp_2 _13265_ (.CLK(clk),
    .D(_01895_),
    .Q(\data_array.data0[11][38] ));
 sky130_fd_sc_hd__dfxtp_2 _13266_ (.CLK(clk),
    .D(_01896_),
    .Q(\data_array.data0[11][39] ));
 sky130_fd_sc_hd__dfxtp_2 _13267_ (.CLK(clk),
    .D(_01897_),
    .Q(\data_array.data0[11][40] ));
 sky130_fd_sc_hd__dfxtp_2 _13268_ (.CLK(clk),
    .D(_01898_),
    .Q(\data_array.data0[11][41] ));
 sky130_fd_sc_hd__dfxtp_2 _13269_ (.CLK(clk),
    .D(_01899_),
    .Q(\data_array.data0[11][42] ));
 sky130_fd_sc_hd__dfxtp_2 _13270_ (.CLK(clk),
    .D(_01900_),
    .Q(\data_array.data0[11][43] ));
 sky130_fd_sc_hd__dfxtp_2 _13271_ (.CLK(clk),
    .D(_01901_),
    .Q(\data_array.data0[11][44] ));
 sky130_fd_sc_hd__dfxtp_2 _13272_ (.CLK(clk),
    .D(_01902_),
    .Q(\data_array.data0[11][45] ));
 sky130_fd_sc_hd__dfxtp_2 _13273_ (.CLK(clk),
    .D(_01903_),
    .Q(\data_array.data0[11][46] ));
 sky130_fd_sc_hd__dfxtp_2 _13274_ (.CLK(clk),
    .D(_01904_),
    .Q(\data_array.data0[11][47] ));
 sky130_fd_sc_hd__dfxtp_2 _13275_ (.CLK(clk),
    .D(_01905_),
    .Q(\data_array.data0[11][48] ));
 sky130_fd_sc_hd__dfxtp_2 _13276_ (.CLK(clk),
    .D(_01906_),
    .Q(\data_array.data0[11][49] ));
 sky130_fd_sc_hd__dfxtp_2 _13277_ (.CLK(clk),
    .D(_01907_),
    .Q(\data_array.data0[11][50] ));
 sky130_fd_sc_hd__dfxtp_2 _13278_ (.CLK(clk),
    .D(_01908_),
    .Q(\data_array.data0[11][51] ));
 sky130_fd_sc_hd__dfxtp_2 _13279_ (.CLK(clk),
    .D(_01909_),
    .Q(\data_array.data0[11][52] ));
 sky130_fd_sc_hd__dfxtp_2 _13280_ (.CLK(clk),
    .D(_01910_),
    .Q(\data_array.data0[11][53] ));
 sky130_fd_sc_hd__dfxtp_2 _13281_ (.CLK(clk),
    .D(_01911_),
    .Q(\data_array.data0[11][54] ));
 sky130_fd_sc_hd__dfxtp_2 _13282_ (.CLK(clk),
    .D(_01912_),
    .Q(\data_array.data0[11][55] ));
 sky130_fd_sc_hd__dfxtp_2 _13283_ (.CLK(clk),
    .D(_01913_),
    .Q(\data_array.data0[11][56] ));
 sky130_fd_sc_hd__dfxtp_2 _13284_ (.CLK(clk),
    .D(_01914_),
    .Q(\data_array.data0[11][57] ));
 sky130_fd_sc_hd__dfxtp_2 _13285_ (.CLK(clk),
    .D(_01915_),
    .Q(\data_array.data0[11][58] ));
 sky130_fd_sc_hd__dfxtp_2 _13286_ (.CLK(clk),
    .D(_01916_),
    .Q(\data_array.data0[11][59] ));
 sky130_fd_sc_hd__dfxtp_2 _13287_ (.CLK(clk),
    .D(_01917_),
    .Q(\data_array.data0[11][60] ));
 sky130_fd_sc_hd__dfxtp_2 _13288_ (.CLK(clk),
    .D(_01918_),
    .Q(\data_array.data0[11][61] ));
 sky130_fd_sc_hd__dfxtp_2 _13289_ (.CLK(clk),
    .D(_01919_),
    .Q(\data_array.data0[11][62] ));
 sky130_fd_sc_hd__dfxtp_2 _13290_ (.CLK(clk),
    .D(_01920_),
    .Q(\data_array.data0[11][63] ));
 sky130_fd_sc_hd__dfxtp_2 _13291_ (.CLK(clk),
    .D(_01921_),
    .Q(\data_array.data0[10][0] ));
 sky130_fd_sc_hd__dfxtp_2 _13292_ (.CLK(clk),
    .D(_01922_),
    .Q(\data_array.data0[10][1] ));
 sky130_fd_sc_hd__dfxtp_2 _13293_ (.CLK(clk),
    .D(_01923_),
    .Q(\data_array.data0[10][2] ));
 sky130_fd_sc_hd__dfxtp_2 _13294_ (.CLK(clk),
    .D(_01924_),
    .Q(\data_array.data0[10][3] ));
 sky130_fd_sc_hd__dfxtp_2 _13295_ (.CLK(clk),
    .D(_01925_),
    .Q(\data_array.data0[10][4] ));
 sky130_fd_sc_hd__dfxtp_2 _13296_ (.CLK(clk),
    .D(_01926_),
    .Q(\data_array.data0[10][5] ));
 sky130_fd_sc_hd__dfxtp_2 _13297_ (.CLK(clk),
    .D(_01927_),
    .Q(\data_array.data0[10][6] ));
 sky130_fd_sc_hd__dfxtp_2 _13298_ (.CLK(clk),
    .D(_01928_),
    .Q(\data_array.data0[10][7] ));
 sky130_fd_sc_hd__dfxtp_2 _13299_ (.CLK(clk),
    .D(_01929_),
    .Q(\data_array.data0[10][8] ));
 sky130_fd_sc_hd__dfxtp_2 _13300_ (.CLK(clk),
    .D(_01930_),
    .Q(\data_array.data0[10][9] ));
 sky130_fd_sc_hd__dfxtp_2 _13301_ (.CLK(clk),
    .D(_01931_),
    .Q(\data_array.data0[10][10] ));
 sky130_fd_sc_hd__dfxtp_2 _13302_ (.CLK(clk),
    .D(_01932_),
    .Q(\data_array.data0[10][11] ));
 sky130_fd_sc_hd__dfxtp_2 _13303_ (.CLK(clk),
    .D(_01933_),
    .Q(\data_array.data0[10][12] ));
 sky130_fd_sc_hd__dfxtp_2 _13304_ (.CLK(clk),
    .D(_01934_),
    .Q(\data_array.data0[10][13] ));
 sky130_fd_sc_hd__dfxtp_2 _13305_ (.CLK(clk),
    .D(_01935_),
    .Q(\data_array.data0[10][14] ));
 sky130_fd_sc_hd__dfxtp_2 _13306_ (.CLK(clk),
    .D(_01936_),
    .Q(\data_array.data0[10][15] ));
 sky130_fd_sc_hd__dfxtp_2 _13307_ (.CLK(clk),
    .D(_01937_),
    .Q(\data_array.data0[10][16] ));
 sky130_fd_sc_hd__dfxtp_2 _13308_ (.CLK(clk),
    .D(_01938_),
    .Q(\data_array.data0[10][17] ));
 sky130_fd_sc_hd__dfxtp_2 _13309_ (.CLK(clk),
    .D(_01939_),
    .Q(\data_array.data0[10][18] ));
 sky130_fd_sc_hd__dfxtp_2 _13310_ (.CLK(clk),
    .D(_01940_),
    .Q(\data_array.data0[10][19] ));
 sky130_fd_sc_hd__dfxtp_2 _13311_ (.CLK(clk),
    .D(_01941_),
    .Q(\data_array.data0[10][20] ));
 sky130_fd_sc_hd__dfxtp_2 _13312_ (.CLK(clk),
    .D(_01942_),
    .Q(\data_array.data0[10][21] ));
 sky130_fd_sc_hd__dfxtp_2 _13313_ (.CLK(clk),
    .D(_01943_),
    .Q(\data_array.data0[10][22] ));
 sky130_fd_sc_hd__dfxtp_2 _13314_ (.CLK(clk),
    .D(_01944_),
    .Q(\data_array.data0[10][23] ));
 sky130_fd_sc_hd__dfxtp_2 _13315_ (.CLK(clk),
    .D(_01945_),
    .Q(\data_array.data0[10][24] ));
 sky130_fd_sc_hd__dfxtp_2 _13316_ (.CLK(clk),
    .D(_01946_),
    .Q(\data_array.data0[10][25] ));
 sky130_fd_sc_hd__dfxtp_2 _13317_ (.CLK(clk),
    .D(_01947_),
    .Q(\data_array.data0[10][26] ));
 sky130_fd_sc_hd__dfxtp_2 _13318_ (.CLK(clk),
    .D(_01948_),
    .Q(\data_array.data0[10][27] ));
 sky130_fd_sc_hd__dfxtp_2 _13319_ (.CLK(clk),
    .D(_01949_),
    .Q(\data_array.data0[10][28] ));
 sky130_fd_sc_hd__dfxtp_2 _13320_ (.CLK(clk),
    .D(_01950_),
    .Q(\data_array.data0[10][29] ));
 sky130_fd_sc_hd__dfxtp_2 _13321_ (.CLK(clk),
    .D(_01951_),
    .Q(\data_array.data0[10][30] ));
 sky130_fd_sc_hd__dfxtp_2 _13322_ (.CLK(clk),
    .D(_01952_),
    .Q(\data_array.data0[10][31] ));
 sky130_fd_sc_hd__dfxtp_2 _13323_ (.CLK(clk),
    .D(_01953_),
    .Q(\data_array.data0[10][32] ));
 sky130_fd_sc_hd__dfxtp_2 _13324_ (.CLK(clk),
    .D(_01954_),
    .Q(\data_array.data0[10][33] ));
 sky130_fd_sc_hd__dfxtp_2 _13325_ (.CLK(clk),
    .D(_01955_),
    .Q(\data_array.data0[10][34] ));
 sky130_fd_sc_hd__dfxtp_2 _13326_ (.CLK(clk),
    .D(_01956_),
    .Q(\data_array.data0[10][35] ));
 sky130_fd_sc_hd__dfxtp_2 _13327_ (.CLK(clk),
    .D(_01957_),
    .Q(\data_array.data0[10][36] ));
 sky130_fd_sc_hd__dfxtp_2 _13328_ (.CLK(clk),
    .D(_01958_),
    .Q(\data_array.data0[10][37] ));
 sky130_fd_sc_hd__dfxtp_2 _13329_ (.CLK(clk),
    .D(_01959_),
    .Q(\data_array.data0[10][38] ));
 sky130_fd_sc_hd__dfxtp_2 _13330_ (.CLK(clk),
    .D(_01960_),
    .Q(\data_array.data0[10][39] ));
 sky130_fd_sc_hd__dfxtp_2 _13331_ (.CLK(clk),
    .D(_01961_),
    .Q(\data_array.data0[10][40] ));
 sky130_fd_sc_hd__dfxtp_2 _13332_ (.CLK(clk),
    .D(_01962_),
    .Q(\data_array.data0[10][41] ));
 sky130_fd_sc_hd__dfxtp_2 _13333_ (.CLK(clk),
    .D(_01963_),
    .Q(\data_array.data0[10][42] ));
 sky130_fd_sc_hd__dfxtp_2 _13334_ (.CLK(clk),
    .D(_01964_),
    .Q(\data_array.data0[10][43] ));
 sky130_fd_sc_hd__dfxtp_2 _13335_ (.CLK(clk),
    .D(_01965_),
    .Q(\data_array.data0[10][44] ));
 sky130_fd_sc_hd__dfxtp_2 _13336_ (.CLK(clk),
    .D(_01966_),
    .Q(\data_array.data0[10][45] ));
 sky130_fd_sc_hd__dfxtp_2 _13337_ (.CLK(clk),
    .D(_01967_),
    .Q(\data_array.data0[10][46] ));
 sky130_fd_sc_hd__dfxtp_2 _13338_ (.CLK(clk),
    .D(_01968_),
    .Q(\data_array.data0[10][47] ));
 sky130_fd_sc_hd__dfxtp_2 _13339_ (.CLK(clk),
    .D(_01969_),
    .Q(\data_array.data0[10][48] ));
 sky130_fd_sc_hd__dfxtp_2 _13340_ (.CLK(clk),
    .D(_01970_),
    .Q(\data_array.data0[10][49] ));
 sky130_fd_sc_hd__dfxtp_2 _13341_ (.CLK(clk),
    .D(_01971_),
    .Q(\data_array.data0[10][50] ));
 sky130_fd_sc_hd__dfxtp_2 _13342_ (.CLK(clk),
    .D(_01972_),
    .Q(\data_array.data0[10][51] ));
 sky130_fd_sc_hd__dfxtp_2 _13343_ (.CLK(clk),
    .D(_01973_),
    .Q(\data_array.data0[10][52] ));
 sky130_fd_sc_hd__dfxtp_2 _13344_ (.CLK(clk),
    .D(_01974_),
    .Q(\data_array.data0[10][53] ));
 sky130_fd_sc_hd__dfxtp_2 _13345_ (.CLK(clk),
    .D(_01975_),
    .Q(\data_array.data0[10][54] ));
 sky130_fd_sc_hd__dfxtp_2 _13346_ (.CLK(clk),
    .D(_01976_),
    .Q(\data_array.data0[10][55] ));
 sky130_fd_sc_hd__dfxtp_2 _13347_ (.CLK(clk),
    .D(_01977_),
    .Q(\data_array.data0[10][56] ));
 sky130_fd_sc_hd__dfxtp_2 _13348_ (.CLK(clk),
    .D(_01978_),
    .Q(\data_array.data0[10][57] ));
 sky130_fd_sc_hd__dfxtp_2 _13349_ (.CLK(clk),
    .D(_01979_),
    .Q(\data_array.data0[10][58] ));
 sky130_fd_sc_hd__dfxtp_2 _13350_ (.CLK(clk),
    .D(_01980_),
    .Q(\data_array.data0[10][59] ));
 sky130_fd_sc_hd__dfxtp_2 _13351_ (.CLK(clk),
    .D(_01981_),
    .Q(\data_array.data0[10][60] ));
 sky130_fd_sc_hd__dfxtp_2 _13352_ (.CLK(clk),
    .D(_01982_),
    .Q(\data_array.data0[10][61] ));
 sky130_fd_sc_hd__dfxtp_2 _13353_ (.CLK(clk),
    .D(_01983_),
    .Q(\data_array.data0[10][62] ));
 sky130_fd_sc_hd__dfxtp_2 _13354_ (.CLK(clk),
    .D(_01984_),
    .Q(\data_array.data0[10][63] ));
 sky130_fd_sc_hd__dfxtp_2 _13355_ (.CLK(clk),
    .D(_01985_),
    .Q(\tag_array.tag0[2][0] ));
 sky130_fd_sc_hd__dfxtp_2 _13356_ (.CLK(clk),
    .D(_01986_),
    .Q(\tag_array.tag0[2][1] ));
 sky130_fd_sc_hd__dfxtp_2 _13357_ (.CLK(clk),
    .D(_01987_),
    .Q(\tag_array.tag0[2][2] ));
 sky130_fd_sc_hd__dfxtp_2 _13358_ (.CLK(clk),
    .D(_01988_),
    .Q(\tag_array.tag0[2][3] ));
 sky130_fd_sc_hd__dfxtp_2 _13359_ (.CLK(clk),
    .D(_01989_),
    .Q(\tag_array.tag0[2][4] ));
 sky130_fd_sc_hd__dfxtp_2 _13360_ (.CLK(clk),
    .D(_01990_),
    .Q(\tag_array.tag0[2][5] ));
 sky130_fd_sc_hd__dfxtp_2 _13361_ (.CLK(clk),
    .D(_01991_),
    .Q(\tag_array.tag0[2][6] ));
 sky130_fd_sc_hd__dfxtp_2 _13362_ (.CLK(clk),
    .D(_01992_),
    .Q(\tag_array.tag0[2][7] ));
 sky130_fd_sc_hd__dfxtp_2 _13363_ (.CLK(clk),
    .D(_01993_),
    .Q(\tag_array.tag0[2][8] ));
 sky130_fd_sc_hd__dfxtp_2 _13364_ (.CLK(clk),
    .D(_01994_),
    .Q(\tag_array.tag0[2][9] ));
 sky130_fd_sc_hd__dfxtp_2 _13365_ (.CLK(clk),
    .D(_01995_),
    .Q(\tag_array.tag0[2][10] ));
 sky130_fd_sc_hd__dfxtp_2 _13366_ (.CLK(clk),
    .D(_01996_),
    .Q(\tag_array.tag0[2][11] ));
 sky130_fd_sc_hd__dfxtp_2 _13367_ (.CLK(clk),
    .D(_01997_),
    .Q(\tag_array.tag0[2][12] ));
 sky130_fd_sc_hd__dfxtp_2 _13368_ (.CLK(clk),
    .D(_01998_),
    .Q(\tag_array.tag0[2][13] ));
 sky130_fd_sc_hd__dfxtp_2 _13369_ (.CLK(clk),
    .D(_01999_),
    .Q(\tag_array.tag0[2][14] ));
 sky130_fd_sc_hd__dfxtp_2 _13370_ (.CLK(clk),
    .D(_02000_),
    .Q(\tag_array.tag0[2][15] ));
 sky130_fd_sc_hd__dfxtp_2 _13371_ (.CLK(clk),
    .D(_02001_),
    .Q(\tag_array.tag0[2][16] ));
 sky130_fd_sc_hd__dfxtp_2 _13372_ (.CLK(clk),
    .D(_02002_),
    .Q(\tag_array.tag0[2][17] ));
 sky130_fd_sc_hd__dfxtp_2 _13373_ (.CLK(clk),
    .D(_02003_),
    .Q(\tag_array.tag0[2][18] ));
 sky130_fd_sc_hd__dfxtp_2 _13374_ (.CLK(clk),
    .D(_02004_),
    .Q(\tag_array.tag0[2][19] ));
 sky130_fd_sc_hd__dfxtp_2 _13375_ (.CLK(clk),
    .D(_02005_),
    .Q(\tag_array.tag0[2][20] ));
 sky130_fd_sc_hd__dfxtp_2 _13376_ (.CLK(clk),
    .D(_02006_),
    .Q(\tag_array.tag0[2][21] ));
 sky130_fd_sc_hd__dfxtp_2 _13377_ (.CLK(clk),
    .D(_02007_),
    .Q(\tag_array.tag0[2][22] ));
 sky130_fd_sc_hd__dfxtp_2 _13378_ (.CLK(clk),
    .D(_02008_),
    .Q(\tag_array.tag0[2][23] ));
 sky130_fd_sc_hd__dfxtp_2 _13379_ (.CLK(clk),
    .D(_02009_),
    .Q(\tag_array.tag0[2][24] ));
 sky130_fd_sc_hd__dfxtp_2 _13380_ (.CLK(clk),
    .D(_02010_),
    .Q(\data_array.data1[8][0] ));
 sky130_fd_sc_hd__dfxtp_2 _13381_ (.CLK(clk),
    .D(_02011_),
    .Q(\data_array.data1[8][1] ));
 sky130_fd_sc_hd__dfxtp_2 _13382_ (.CLK(clk),
    .D(_02012_),
    .Q(\data_array.data1[8][2] ));
 sky130_fd_sc_hd__dfxtp_2 _13383_ (.CLK(clk),
    .D(_02013_),
    .Q(\data_array.data1[8][3] ));
 sky130_fd_sc_hd__dfxtp_2 _13384_ (.CLK(clk),
    .D(_02014_),
    .Q(\data_array.data1[8][4] ));
 sky130_fd_sc_hd__dfxtp_2 _13385_ (.CLK(clk),
    .D(_02015_),
    .Q(\data_array.data1[8][5] ));
 sky130_fd_sc_hd__dfxtp_2 _13386_ (.CLK(clk),
    .D(_02016_),
    .Q(\data_array.data1[8][6] ));
 sky130_fd_sc_hd__dfxtp_2 _13387_ (.CLK(clk),
    .D(_02017_),
    .Q(\data_array.data1[8][7] ));
 sky130_fd_sc_hd__dfxtp_2 _13388_ (.CLK(clk),
    .D(_02018_),
    .Q(\data_array.data1[8][8] ));
 sky130_fd_sc_hd__dfxtp_2 _13389_ (.CLK(clk),
    .D(_02019_),
    .Q(\data_array.data1[8][9] ));
 sky130_fd_sc_hd__dfxtp_2 _13390_ (.CLK(clk),
    .D(_02020_),
    .Q(\data_array.data1[8][10] ));
 sky130_fd_sc_hd__dfxtp_2 _13391_ (.CLK(clk),
    .D(_02021_),
    .Q(\data_array.data1[8][11] ));
 sky130_fd_sc_hd__dfxtp_2 _13392_ (.CLK(clk),
    .D(_02022_),
    .Q(\data_array.data1[8][12] ));
 sky130_fd_sc_hd__dfxtp_2 _13393_ (.CLK(clk),
    .D(_02023_),
    .Q(\data_array.data1[8][13] ));
 sky130_fd_sc_hd__dfxtp_2 _13394_ (.CLK(clk),
    .D(_02024_),
    .Q(\data_array.data1[8][14] ));
 sky130_fd_sc_hd__dfxtp_2 _13395_ (.CLK(clk),
    .D(_02025_),
    .Q(\data_array.data1[8][15] ));
 sky130_fd_sc_hd__dfxtp_2 _13396_ (.CLK(clk),
    .D(_02026_),
    .Q(\data_array.data1[8][16] ));
 sky130_fd_sc_hd__dfxtp_2 _13397_ (.CLK(clk),
    .D(_02027_),
    .Q(\data_array.data1[8][17] ));
 sky130_fd_sc_hd__dfxtp_2 _13398_ (.CLK(clk),
    .D(_02028_),
    .Q(\data_array.data1[8][18] ));
 sky130_fd_sc_hd__dfxtp_2 _13399_ (.CLK(clk),
    .D(_02029_),
    .Q(\data_array.data1[8][19] ));
 sky130_fd_sc_hd__dfxtp_2 _13400_ (.CLK(clk),
    .D(_02030_),
    .Q(\data_array.data1[8][20] ));
 sky130_fd_sc_hd__dfxtp_2 _13401_ (.CLK(clk),
    .D(_02031_),
    .Q(\data_array.data1[8][21] ));
 sky130_fd_sc_hd__dfxtp_2 _13402_ (.CLK(clk),
    .D(_02032_),
    .Q(\data_array.data1[8][22] ));
 sky130_fd_sc_hd__dfxtp_2 _13403_ (.CLK(clk),
    .D(_02033_),
    .Q(\data_array.data1[8][23] ));
 sky130_fd_sc_hd__dfxtp_2 _13404_ (.CLK(clk),
    .D(_02034_),
    .Q(\data_array.data1[8][24] ));
 sky130_fd_sc_hd__dfxtp_2 _13405_ (.CLK(clk),
    .D(_02035_),
    .Q(\data_array.data1[8][25] ));
 sky130_fd_sc_hd__dfxtp_2 _13406_ (.CLK(clk),
    .D(_02036_),
    .Q(\data_array.data1[8][26] ));
 sky130_fd_sc_hd__dfxtp_2 _13407_ (.CLK(clk),
    .D(_02037_),
    .Q(\data_array.data1[8][27] ));
 sky130_fd_sc_hd__dfxtp_2 _13408_ (.CLK(clk),
    .D(_02038_),
    .Q(\data_array.data1[8][28] ));
 sky130_fd_sc_hd__dfxtp_2 _13409_ (.CLK(clk),
    .D(_02039_),
    .Q(\data_array.data1[8][29] ));
 sky130_fd_sc_hd__dfxtp_2 _13410_ (.CLK(clk),
    .D(_02040_),
    .Q(\data_array.data1[8][30] ));
 sky130_fd_sc_hd__dfxtp_2 _13411_ (.CLK(clk),
    .D(_02041_),
    .Q(\data_array.data1[8][31] ));
 sky130_fd_sc_hd__dfxtp_2 _13412_ (.CLK(clk),
    .D(_02042_),
    .Q(\data_array.data1[8][32] ));
 sky130_fd_sc_hd__dfxtp_2 _13413_ (.CLK(clk),
    .D(_02043_),
    .Q(\data_array.data1[8][33] ));
 sky130_fd_sc_hd__dfxtp_2 _13414_ (.CLK(clk),
    .D(_02044_),
    .Q(\data_array.data1[8][34] ));
 sky130_fd_sc_hd__dfxtp_2 _13415_ (.CLK(clk),
    .D(_02045_),
    .Q(\data_array.data1[8][35] ));
 sky130_fd_sc_hd__dfxtp_2 _13416_ (.CLK(clk),
    .D(_02046_),
    .Q(\data_array.data1[8][36] ));
 sky130_fd_sc_hd__dfxtp_2 _13417_ (.CLK(clk),
    .D(_02047_),
    .Q(\data_array.data1[8][37] ));
 sky130_fd_sc_hd__dfxtp_2 _13418_ (.CLK(clk),
    .D(_02048_),
    .Q(\data_array.data1[8][38] ));
 sky130_fd_sc_hd__dfxtp_2 _13419_ (.CLK(clk),
    .D(_02049_),
    .Q(\data_array.data1[8][39] ));
 sky130_fd_sc_hd__dfxtp_2 _13420_ (.CLK(clk),
    .D(_02050_),
    .Q(\data_array.data1[8][40] ));
 sky130_fd_sc_hd__dfxtp_2 _13421_ (.CLK(clk),
    .D(_02051_),
    .Q(\data_array.data1[8][41] ));
 sky130_fd_sc_hd__dfxtp_2 _13422_ (.CLK(clk),
    .D(_02052_),
    .Q(\data_array.data1[8][42] ));
 sky130_fd_sc_hd__dfxtp_2 _13423_ (.CLK(clk),
    .D(_02053_),
    .Q(\data_array.data1[8][43] ));
 sky130_fd_sc_hd__dfxtp_2 _13424_ (.CLK(clk),
    .D(_02054_),
    .Q(\data_array.data1[8][44] ));
 sky130_fd_sc_hd__dfxtp_2 _13425_ (.CLK(clk),
    .D(_02055_),
    .Q(\data_array.data1[8][45] ));
 sky130_fd_sc_hd__dfxtp_2 _13426_ (.CLK(clk),
    .D(_02056_),
    .Q(\data_array.data1[8][46] ));
 sky130_fd_sc_hd__dfxtp_2 _13427_ (.CLK(clk),
    .D(_02057_),
    .Q(\data_array.data1[8][47] ));
 sky130_fd_sc_hd__dfxtp_2 _13428_ (.CLK(clk),
    .D(_02058_),
    .Q(\data_array.data1[8][48] ));
 sky130_fd_sc_hd__dfxtp_2 _13429_ (.CLK(clk),
    .D(_02059_),
    .Q(\data_array.data1[8][49] ));
 sky130_fd_sc_hd__dfxtp_2 _13430_ (.CLK(clk),
    .D(_02060_),
    .Q(\data_array.data1[8][50] ));
 sky130_fd_sc_hd__dfxtp_2 _13431_ (.CLK(clk),
    .D(_02061_),
    .Q(\data_array.data1[8][51] ));
 sky130_fd_sc_hd__dfxtp_2 _13432_ (.CLK(clk),
    .D(_02062_),
    .Q(\data_array.data1[8][52] ));
 sky130_fd_sc_hd__dfxtp_2 _13433_ (.CLK(clk),
    .D(_02063_),
    .Q(\data_array.data1[8][53] ));
 sky130_fd_sc_hd__dfxtp_2 _13434_ (.CLK(clk),
    .D(_02064_),
    .Q(\data_array.data1[8][54] ));
 sky130_fd_sc_hd__dfxtp_2 _13435_ (.CLK(clk),
    .D(_02065_),
    .Q(\data_array.data1[8][55] ));
 sky130_fd_sc_hd__dfxtp_2 _13436_ (.CLK(clk),
    .D(_02066_),
    .Q(\data_array.data1[8][56] ));
 sky130_fd_sc_hd__dfxtp_2 _13437_ (.CLK(clk),
    .D(_02067_),
    .Q(\data_array.data1[8][57] ));
 sky130_fd_sc_hd__dfxtp_2 _13438_ (.CLK(clk),
    .D(_02068_),
    .Q(\data_array.data1[8][58] ));
 sky130_fd_sc_hd__dfxtp_2 _13439_ (.CLK(clk),
    .D(_02069_),
    .Q(\data_array.data1[8][59] ));
 sky130_fd_sc_hd__dfxtp_2 _13440_ (.CLK(clk),
    .D(_02070_),
    .Q(\data_array.data1[8][60] ));
 sky130_fd_sc_hd__dfxtp_2 _13441_ (.CLK(clk),
    .D(_02071_),
    .Q(\data_array.data1[8][61] ));
 sky130_fd_sc_hd__dfxtp_2 _13442_ (.CLK(clk),
    .D(_02072_),
    .Q(\data_array.data1[8][62] ));
 sky130_fd_sc_hd__dfxtp_2 _13443_ (.CLK(clk),
    .D(_02073_),
    .Q(\data_array.data1[8][63] ));
 sky130_fd_sc_hd__dfxtp_2 _13444_ (.CLK(clk),
    .D(_02074_),
    .Q(\tag_array.tag0[1][0] ));
 sky130_fd_sc_hd__dfxtp_2 _13445_ (.CLK(clk),
    .D(_02075_),
    .Q(\tag_array.tag0[1][1] ));
 sky130_fd_sc_hd__dfxtp_2 _13446_ (.CLK(clk),
    .D(_02076_),
    .Q(\tag_array.tag0[1][2] ));
 sky130_fd_sc_hd__dfxtp_2 _13447_ (.CLK(clk),
    .D(_02077_),
    .Q(\tag_array.tag0[1][3] ));
 sky130_fd_sc_hd__dfxtp_2 _13448_ (.CLK(clk),
    .D(_02078_),
    .Q(\tag_array.tag0[1][4] ));
 sky130_fd_sc_hd__dfxtp_2 _13449_ (.CLK(clk),
    .D(_02079_),
    .Q(\tag_array.tag0[1][5] ));
 sky130_fd_sc_hd__dfxtp_2 _13450_ (.CLK(clk),
    .D(_02080_),
    .Q(\tag_array.tag0[1][6] ));
 sky130_fd_sc_hd__dfxtp_2 _13451_ (.CLK(clk),
    .D(_02081_),
    .Q(\tag_array.tag0[1][7] ));
 sky130_fd_sc_hd__dfxtp_2 _13452_ (.CLK(clk),
    .D(_02082_),
    .Q(\tag_array.tag0[1][8] ));
 sky130_fd_sc_hd__dfxtp_2 _13453_ (.CLK(clk),
    .D(_02083_),
    .Q(\tag_array.tag0[1][9] ));
 sky130_fd_sc_hd__dfxtp_2 _13454_ (.CLK(clk),
    .D(_02084_),
    .Q(\tag_array.tag0[1][10] ));
 sky130_fd_sc_hd__dfxtp_2 _13455_ (.CLK(clk),
    .D(_02085_),
    .Q(\tag_array.tag0[1][11] ));
 sky130_fd_sc_hd__dfxtp_2 _13456_ (.CLK(clk),
    .D(_02086_),
    .Q(\tag_array.tag0[1][12] ));
 sky130_fd_sc_hd__dfxtp_2 _13457_ (.CLK(clk),
    .D(_02087_),
    .Q(\tag_array.tag0[1][13] ));
 sky130_fd_sc_hd__dfxtp_2 _13458_ (.CLK(clk),
    .D(_02088_),
    .Q(\tag_array.tag0[1][14] ));
 sky130_fd_sc_hd__dfxtp_2 _13459_ (.CLK(clk),
    .D(_02089_),
    .Q(\tag_array.tag0[1][15] ));
 sky130_fd_sc_hd__dfxtp_2 _13460_ (.CLK(clk),
    .D(_02090_),
    .Q(\tag_array.tag0[1][16] ));
 sky130_fd_sc_hd__dfxtp_2 _13461_ (.CLK(clk),
    .D(_02091_),
    .Q(\tag_array.tag0[1][17] ));
 sky130_fd_sc_hd__dfxtp_2 _13462_ (.CLK(clk),
    .D(_02092_),
    .Q(\tag_array.tag0[1][18] ));
 sky130_fd_sc_hd__dfxtp_2 _13463_ (.CLK(clk),
    .D(_02093_),
    .Q(\tag_array.tag0[1][19] ));
 sky130_fd_sc_hd__dfxtp_2 _13464_ (.CLK(clk),
    .D(_02094_),
    .Q(\tag_array.tag0[1][20] ));
 sky130_fd_sc_hd__dfxtp_2 _13465_ (.CLK(clk),
    .D(_02095_),
    .Q(\tag_array.tag0[1][21] ));
 sky130_fd_sc_hd__dfxtp_2 _13466_ (.CLK(clk),
    .D(_02096_),
    .Q(\tag_array.tag0[1][22] ));
 sky130_fd_sc_hd__dfxtp_2 _13467_ (.CLK(clk),
    .D(_02097_),
    .Q(\tag_array.tag0[1][23] ));
 sky130_fd_sc_hd__dfxtp_2 _13468_ (.CLK(clk),
    .D(_02098_),
    .Q(\tag_array.tag0[1][24] ));
 sky130_fd_sc_hd__dfxtp_2 _13469_ (.CLK(clk),
    .D(_02099_),
    .Q(\tag_array.tag0[15][0] ));
 sky130_fd_sc_hd__dfxtp_2 _13470_ (.CLK(clk),
    .D(_02100_),
    .Q(\tag_array.tag0[15][1] ));
 sky130_fd_sc_hd__dfxtp_2 _13471_ (.CLK(clk),
    .D(_02101_),
    .Q(\tag_array.tag0[15][2] ));
 sky130_fd_sc_hd__dfxtp_2 _13472_ (.CLK(clk),
    .D(_02102_),
    .Q(\tag_array.tag0[15][3] ));
 sky130_fd_sc_hd__dfxtp_2 _13473_ (.CLK(clk),
    .D(_02103_),
    .Q(\tag_array.tag0[15][4] ));
 sky130_fd_sc_hd__dfxtp_2 _13474_ (.CLK(clk),
    .D(_02104_),
    .Q(\tag_array.tag0[15][5] ));
 sky130_fd_sc_hd__dfxtp_2 _13475_ (.CLK(clk),
    .D(_02105_),
    .Q(\tag_array.tag0[15][6] ));
 sky130_fd_sc_hd__dfxtp_2 _13476_ (.CLK(clk),
    .D(_02106_),
    .Q(\tag_array.tag0[15][7] ));
 sky130_fd_sc_hd__dfxtp_2 _13477_ (.CLK(clk),
    .D(_02107_),
    .Q(\tag_array.tag0[15][8] ));
 sky130_fd_sc_hd__dfxtp_2 _13478_ (.CLK(clk),
    .D(_02108_),
    .Q(\tag_array.tag0[15][9] ));
 sky130_fd_sc_hd__dfxtp_2 _13479_ (.CLK(clk),
    .D(_02109_),
    .Q(\tag_array.tag0[15][10] ));
 sky130_fd_sc_hd__dfxtp_2 _13480_ (.CLK(clk),
    .D(_02110_),
    .Q(\tag_array.tag0[15][11] ));
 sky130_fd_sc_hd__dfxtp_2 _13481_ (.CLK(clk),
    .D(_02111_),
    .Q(\tag_array.tag0[15][12] ));
 sky130_fd_sc_hd__dfxtp_2 _13482_ (.CLK(clk),
    .D(_02112_),
    .Q(\tag_array.tag0[15][13] ));
 sky130_fd_sc_hd__dfxtp_2 _13483_ (.CLK(clk),
    .D(_02113_),
    .Q(\tag_array.tag0[15][14] ));
 sky130_fd_sc_hd__dfxtp_2 _13484_ (.CLK(clk),
    .D(_02114_),
    .Q(\tag_array.tag0[15][15] ));
 sky130_fd_sc_hd__dfxtp_2 _13485_ (.CLK(clk),
    .D(_02115_),
    .Q(\tag_array.tag0[15][16] ));
 sky130_fd_sc_hd__dfxtp_2 _13486_ (.CLK(clk),
    .D(_02116_),
    .Q(\tag_array.tag0[15][17] ));
 sky130_fd_sc_hd__dfxtp_2 _13487_ (.CLK(clk),
    .D(_02117_),
    .Q(\tag_array.tag0[15][18] ));
 sky130_fd_sc_hd__dfxtp_2 _13488_ (.CLK(clk),
    .D(_02118_),
    .Q(\tag_array.tag0[15][19] ));
 sky130_fd_sc_hd__dfxtp_2 _13489_ (.CLK(clk),
    .D(_02119_),
    .Q(\tag_array.tag0[15][20] ));
 sky130_fd_sc_hd__dfxtp_2 _13490_ (.CLK(clk),
    .D(_02120_),
    .Q(\tag_array.tag0[15][21] ));
 sky130_fd_sc_hd__dfxtp_2 _13491_ (.CLK(clk),
    .D(_02121_),
    .Q(\tag_array.tag0[15][22] ));
 sky130_fd_sc_hd__dfxtp_2 _13492_ (.CLK(clk),
    .D(_02122_),
    .Q(\tag_array.tag0[15][23] ));
 sky130_fd_sc_hd__dfxtp_2 _13493_ (.CLK(clk),
    .D(_02123_),
    .Q(\tag_array.tag0[15][24] ));
 sky130_fd_sc_hd__dfxtp_2 _13494_ (.CLK(clk),
    .D(_02124_),
    .Q(\tag_array.dirty1[9] ));
 sky130_fd_sc_hd__dfxtp_2 _13495_ (.CLK(clk),
    .D(_00130_),
    .Q(dirty_way1));
 sky130_fd_sc_hd__dfxtp_2 _13496_ (.CLK(clk),
    .D(_02125_),
    .Q(\tag_array.dirty1[14] ));
 sky130_fd_sc_hd__dfxtp_2 _13497_ (.CLK(clk),
    .D(_02126_),
    .Q(\tag_array.dirty1[13] ));
 sky130_fd_sc_hd__dfxtp_2 _13498_ (.CLK(clk),
    .D(_02127_),
    .Q(\tag_array.dirty1[12] ));
 sky130_fd_sc_hd__dfxtp_2 _13499_ (.CLK(clk),
    .D(_02128_),
    .Q(\tag_array.dirty1[11] ));
 sky130_fd_sc_hd__dfxtp_2 _13500_ (.CLK(clk),
    .D(_02129_),
    .Q(\tag_array.dirty1[10] ));
 sky130_fd_sc_hd__dfxtp_2 _13501_ (.CLK(clk),
    .D(_02130_),
    .Q(\tag_array.dirty1[0] ));
 sky130_fd_sc_hd__dfxtp_2 _13502_ (.CLK(clk),
    .D(_02131_),
    .Q(\tag_array.dirty1[8] ));
 sky130_fd_sc_hd__dfxtp_2 _13503_ (.CLK(clk),
    .D(_02132_),
    .Q(\data_array.data1[0][0] ));
 sky130_fd_sc_hd__dfxtp_2 _13504_ (.CLK(clk),
    .D(_02133_),
    .Q(\data_array.data1[0][1] ));
 sky130_fd_sc_hd__dfxtp_2 _13505_ (.CLK(clk),
    .D(_02134_),
    .Q(\data_array.data1[0][2] ));
 sky130_fd_sc_hd__dfxtp_2 _13506_ (.CLK(clk),
    .D(_02135_),
    .Q(\data_array.data1[0][3] ));
 sky130_fd_sc_hd__dfxtp_2 _13507_ (.CLK(clk),
    .D(_02136_),
    .Q(\data_array.data1[0][4] ));
 sky130_fd_sc_hd__dfxtp_2 _13508_ (.CLK(clk),
    .D(_02137_),
    .Q(\data_array.data1[0][5] ));
 sky130_fd_sc_hd__dfxtp_2 _13509_ (.CLK(clk),
    .D(_02138_),
    .Q(\data_array.data1[0][6] ));
 sky130_fd_sc_hd__dfxtp_2 _13510_ (.CLK(clk),
    .D(_02139_),
    .Q(\data_array.data1[0][7] ));
 sky130_fd_sc_hd__dfxtp_2 _13511_ (.CLK(clk),
    .D(_02140_),
    .Q(\data_array.data1[0][8] ));
 sky130_fd_sc_hd__dfxtp_2 _13512_ (.CLK(clk),
    .D(_02141_),
    .Q(\data_array.data1[0][9] ));
 sky130_fd_sc_hd__dfxtp_2 _13513_ (.CLK(clk),
    .D(_02142_),
    .Q(\data_array.data1[0][10] ));
 sky130_fd_sc_hd__dfxtp_2 _13514_ (.CLK(clk),
    .D(_02143_),
    .Q(\data_array.data1[0][11] ));
 sky130_fd_sc_hd__dfxtp_2 _13515_ (.CLK(clk),
    .D(_02144_),
    .Q(\data_array.data1[0][12] ));
 sky130_fd_sc_hd__dfxtp_2 _13516_ (.CLK(clk),
    .D(_02145_),
    .Q(\data_array.data1[0][13] ));
 sky130_fd_sc_hd__dfxtp_2 _13517_ (.CLK(clk),
    .D(_02146_),
    .Q(\data_array.data1[0][14] ));
 sky130_fd_sc_hd__dfxtp_2 _13518_ (.CLK(clk),
    .D(_02147_),
    .Q(\data_array.data1[0][15] ));
 sky130_fd_sc_hd__dfxtp_2 _13519_ (.CLK(clk),
    .D(_02148_),
    .Q(\data_array.data1[0][16] ));
 sky130_fd_sc_hd__dfxtp_2 _13520_ (.CLK(clk),
    .D(_02149_),
    .Q(\data_array.data1[0][17] ));
 sky130_fd_sc_hd__dfxtp_2 _13521_ (.CLK(clk),
    .D(_02150_),
    .Q(\data_array.data1[0][18] ));
 sky130_fd_sc_hd__dfxtp_2 _13522_ (.CLK(clk),
    .D(_02151_),
    .Q(\data_array.data1[0][19] ));
 sky130_fd_sc_hd__dfxtp_2 _13523_ (.CLK(clk),
    .D(_02152_),
    .Q(\data_array.data1[0][20] ));
 sky130_fd_sc_hd__dfxtp_2 _13524_ (.CLK(clk),
    .D(_02153_),
    .Q(\data_array.data1[0][21] ));
 sky130_fd_sc_hd__dfxtp_2 _13525_ (.CLK(clk),
    .D(_02154_),
    .Q(\data_array.data1[0][22] ));
 sky130_fd_sc_hd__dfxtp_2 _13526_ (.CLK(clk),
    .D(_02155_),
    .Q(\data_array.data1[0][23] ));
 sky130_fd_sc_hd__dfxtp_2 _13527_ (.CLK(clk),
    .D(_02156_),
    .Q(\data_array.data1[0][24] ));
 sky130_fd_sc_hd__dfxtp_2 _13528_ (.CLK(clk),
    .D(_02157_),
    .Q(\data_array.data1[0][25] ));
 sky130_fd_sc_hd__dfxtp_2 _13529_ (.CLK(clk),
    .D(_02158_),
    .Q(\data_array.data1[0][26] ));
 sky130_fd_sc_hd__dfxtp_2 _13530_ (.CLK(clk),
    .D(_02159_),
    .Q(\data_array.data1[0][27] ));
 sky130_fd_sc_hd__dfxtp_2 _13531_ (.CLK(clk),
    .D(_02160_),
    .Q(\data_array.data1[0][28] ));
 sky130_fd_sc_hd__dfxtp_2 _13532_ (.CLK(clk),
    .D(_02161_),
    .Q(\data_array.data1[0][29] ));
 sky130_fd_sc_hd__dfxtp_2 _13533_ (.CLK(clk),
    .D(_02162_),
    .Q(\data_array.data1[0][30] ));
 sky130_fd_sc_hd__dfxtp_2 _13534_ (.CLK(clk),
    .D(_02163_),
    .Q(\data_array.data1[0][31] ));
 sky130_fd_sc_hd__dfxtp_2 _13535_ (.CLK(clk),
    .D(_02164_),
    .Q(\data_array.data1[0][32] ));
 sky130_fd_sc_hd__dfxtp_2 _13536_ (.CLK(clk),
    .D(_02165_),
    .Q(\data_array.data1[0][33] ));
 sky130_fd_sc_hd__dfxtp_2 _13537_ (.CLK(clk),
    .D(_02166_),
    .Q(\data_array.data1[0][34] ));
 sky130_fd_sc_hd__dfxtp_2 _13538_ (.CLK(clk),
    .D(_02167_),
    .Q(\data_array.data1[0][35] ));
 sky130_fd_sc_hd__dfxtp_2 _13539_ (.CLK(clk),
    .D(_02168_),
    .Q(\data_array.data1[0][36] ));
 sky130_fd_sc_hd__dfxtp_2 _13540_ (.CLK(clk),
    .D(_02169_),
    .Q(\data_array.data1[0][37] ));
 sky130_fd_sc_hd__dfxtp_2 _13541_ (.CLK(clk),
    .D(_02170_),
    .Q(\data_array.data1[0][38] ));
 sky130_fd_sc_hd__dfxtp_2 _13542_ (.CLK(clk),
    .D(_02171_),
    .Q(\data_array.data1[0][39] ));
 sky130_fd_sc_hd__dfxtp_2 _13543_ (.CLK(clk),
    .D(_02172_),
    .Q(\data_array.data1[0][40] ));
 sky130_fd_sc_hd__dfxtp_2 _13544_ (.CLK(clk),
    .D(_02173_),
    .Q(\data_array.data1[0][41] ));
 sky130_fd_sc_hd__dfxtp_2 _13545_ (.CLK(clk),
    .D(_02174_),
    .Q(\data_array.data1[0][42] ));
 sky130_fd_sc_hd__dfxtp_2 _13546_ (.CLK(clk),
    .D(_02175_),
    .Q(\data_array.data1[0][43] ));
 sky130_fd_sc_hd__dfxtp_2 _13547_ (.CLK(clk),
    .D(_02176_),
    .Q(\data_array.data1[0][44] ));
 sky130_fd_sc_hd__dfxtp_2 _13548_ (.CLK(clk),
    .D(_02177_),
    .Q(\data_array.data1[0][45] ));
 sky130_fd_sc_hd__dfxtp_2 _13549_ (.CLK(clk),
    .D(_02178_),
    .Q(\data_array.data1[0][46] ));
 sky130_fd_sc_hd__dfxtp_2 _13550_ (.CLK(clk),
    .D(_02179_),
    .Q(\data_array.data1[0][47] ));
 sky130_fd_sc_hd__dfxtp_2 _13551_ (.CLK(clk),
    .D(_02180_),
    .Q(\data_array.data1[0][48] ));
 sky130_fd_sc_hd__dfxtp_2 _13552_ (.CLK(clk),
    .D(_02181_),
    .Q(\data_array.data1[0][49] ));
 sky130_fd_sc_hd__dfxtp_2 _13553_ (.CLK(clk),
    .D(_02182_),
    .Q(\data_array.data1[0][50] ));
 sky130_fd_sc_hd__dfxtp_2 _13554_ (.CLK(clk),
    .D(_02183_),
    .Q(\data_array.data1[0][51] ));
 sky130_fd_sc_hd__dfxtp_2 _13555_ (.CLK(clk),
    .D(_02184_),
    .Q(\data_array.data1[0][52] ));
 sky130_fd_sc_hd__dfxtp_2 _13556_ (.CLK(clk),
    .D(_02185_),
    .Q(\data_array.data1[0][53] ));
 sky130_fd_sc_hd__dfxtp_2 _13557_ (.CLK(clk),
    .D(_02186_),
    .Q(\data_array.data1[0][54] ));
 sky130_fd_sc_hd__dfxtp_2 _13558_ (.CLK(clk),
    .D(_02187_),
    .Q(\data_array.data1[0][55] ));
 sky130_fd_sc_hd__dfxtp_2 _13559_ (.CLK(clk),
    .D(_02188_),
    .Q(\data_array.data1[0][56] ));
 sky130_fd_sc_hd__dfxtp_2 _13560_ (.CLK(clk),
    .D(_02189_),
    .Q(\data_array.data1[0][57] ));
 sky130_fd_sc_hd__dfxtp_2 _13561_ (.CLK(clk),
    .D(_02190_),
    .Q(\data_array.data1[0][58] ));
 sky130_fd_sc_hd__dfxtp_2 _13562_ (.CLK(clk),
    .D(_02191_),
    .Q(\data_array.data1[0][59] ));
 sky130_fd_sc_hd__dfxtp_2 _13563_ (.CLK(clk),
    .D(_02192_),
    .Q(\data_array.data1[0][60] ));
 sky130_fd_sc_hd__dfxtp_2 _13564_ (.CLK(clk),
    .D(_02193_),
    .Q(\data_array.data1[0][61] ));
 sky130_fd_sc_hd__dfxtp_2 _13565_ (.CLK(clk),
    .D(_02194_),
    .Q(\data_array.data1[0][62] ));
 sky130_fd_sc_hd__dfxtp_2 _13566_ (.CLK(clk),
    .D(_02195_),
    .Q(\data_array.data1[0][63] ));
 sky130_fd_sc_hd__dfxtp_2 _13567_ (.CLK(clk),
    .D(_02196_),
    .Q(\tag_array.dirty1[7] ));
 sky130_fd_sc_hd__dfxtp_2 _13568_ (.CLK(clk),
    .D(_02197_),
    .Q(\tag_array.dirty1[6] ));
 sky130_fd_sc_hd__dfxtp_2 _13569_ (.CLK(clk),
    .D(_02198_),
    .Q(\tag_array.dirty1[5] ));
 sky130_fd_sc_hd__dfxtp_2 _13570_ (.CLK(clk),
    .D(_02199_),
    .Q(\tag_array.dirty1[4] ));
 sky130_fd_sc_hd__dfxtp_2 _13571_ (.CLK(clk),
    .D(_02200_),
    .Q(\tag_array.dirty1[3] ));
 sky130_fd_sc_hd__dfxtp_2 _13572_ (.CLK(clk),
    .D(_02201_),
    .Q(\tag_array.dirty1[2] ));
 sky130_fd_sc_hd__dfxtp_2 _13573_ (.CLK(clk),
    .D(_02202_),
    .Q(\tag_array.dirty1[1] ));
 sky130_fd_sc_hd__dfxtp_2 _13574_ (.CLK(clk),
    .D(_02203_),
    .Q(\tag_array.dirty1[15] ));
 sky130_fd_sc_hd__dfxtp_2 _13575_ (.CLK(clk),
    .D(_02204_),
    .Q(\data_array.data0[9][0] ));
 sky130_fd_sc_hd__dfxtp_2 _13576_ (.CLK(clk),
    .D(_02205_),
    .Q(\data_array.data0[9][1] ));
 sky130_fd_sc_hd__dfxtp_2 _13577_ (.CLK(clk),
    .D(_02206_),
    .Q(\data_array.data0[9][2] ));
 sky130_fd_sc_hd__dfxtp_2 _13578_ (.CLK(clk),
    .D(_02207_),
    .Q(\data_array.data0[9][3] ));
 sky130_fd_sc_hd__dfxtp_2 _13579_ (.CLK(clk),
    .D(_02208_),
    .Q(\data_array.data0[9][4] ));
 sky130_fd_sc_hd__dfxtp_2 _13580_ (.CLK(clk),
    .D(_02209_),
    .Q(\data_array.data0[9][5] ));
 sky130_fd_sc_hd__dfxtp_2 _13581_ (.CLK(clk),
    .D(_02210_),
    .Q(\data_array.data0[9][6] ));
 sky130_fd_sc_hd__dfxtp_2 _13582_ (.CLK(clk),
    .D(_02211_),
    .Q(\data_array.data0[9][7] ));
 sky130_fd_sc_hd__dfxtp_2 _13583_ (.CLK(clk),
    .D(_02212_),
    .Q(\data_array.data0[9][8] ));
 sky130_fd_sc_hd__dfxtp_2 _13584_ (.CLK(clk),
    .D(_02213_),
    .Q(\data_array.data0[9][9] ));
 sky130_fd_sc_hd__dfxtp_2 _13585_ (.CLK(clk),
    .D(_02214_),
    .Q(\data_array.data0[9][10] ));
 sky130_fd_sc_hd__dfxtp_2 _13586_ (.CLK(clk),
    .D(_02215_),
    .Q(\data_array.data0[9][11] ));
 sky130_fd_sc_hd__dfxtp_2 _13587_ (.CLK(clk),
    .D(_02216_),
    .Q(\data_array.data0[9][12] ));
 sky130_fd_sc_hd__dfxtp_2 _13588_ (.CLK(clk),
    .D(_02217_),
    .Q(\data_array.data0[9][13] ));
 sky130_fd_sc_hd__dfxtp_2 _13589_ (.CLK(clk),
    .D(_02218_),
    .Q(\data_array.data0[9][14] ));
 sky130_fd_sc_hd__dfxtp_2 _13590_ (.CLK(clk),
    .D(_02219_),
    .Q(\data_array.data0[9][15] ));
 sky130_fd_sc_hd__dfxtp_2 _13591_ (.CLK(clk),
    .D(_02220_),
    .Q(\data_array.data0[9][16] ));
 sky130_fd_sc_hd__dfxtp_2 _13592_ (.CLK(clk),
    .D(_02221_),
    .Q(\data_array.data0[9][17] ));
 sky130_fd_sc_hd__dfxtp_2 _13593_ (.CLK(clk),
    .D(_02222_),
    .Q(\data_array.data0[9][18] ));
 sky130_fd_sc_hd__dfxtp_2 _13594_ (.CLK(clk),
    .D(_02223_),
    .Q(\data_array.data0[9][19] ));
 sky130_fd_sc_hd__dfxtp_2 _13595_ (.CLK(clk),
    .D(_02224_),
    .Q(\data_array.data0[9][20] ));
 sky130_fd_sc_hd__dfxtp_2 _13596_ (.CLK(clk),
    .D(_02225_),
    .Q(\data_array.data0[9][21] ));
 sky130_fd_sc_hd__dfxtp_2 _13597_ (.CLK(clk),
    .D(_02226_),
    .Q(\data_array.data0[9][22] ));
 sky130_fd_sc_hd__dfxtp_2 _13598_ (.CLK(clk),
    .D(_02227_),
    .Q(\data_array.data0[9][23] ));
 sky130_fd_sc_hd__dfxtp_2 _13599_ (.CLK(clk),
    .D(_02228_),
    .Q(\data_array.data0[9][24] ));
 sky130_fd_sc_hd__dfxtp_2 _13600_ (.CLK(clk),
    .D(_02229_),
    .Q(\data_array.data0[9][25] ));
 sky130_fd_sc_hd__dfxtp_2 _13601_ (.CLK(clk),
    .D(_02230_),
    .Q(\data_array.data0[9][26] ));
 sky130_fd_sc_hd__dfxtp_2 _13602_ (.CLK(clk),
    .D(_02231_),
    .Q(\data_array.data0[9][27] ));
 sky130_fd_sc_hd__dfxtp_2 _13603_ (.CLK(clk),
    .D(_02232_),
    .Q(\data_array.data0[9][28] ));
 sky130_fd_sc_hd__dfxtp_2 _13604_ (.CLK(clk),
    .D(_02233_),
    .Q(\data_array.data0[9][29] ));
 sky130_fd_sc_hd__dfxtp_2 _13605_ (.CLK(clk),
    .D(_02234_),
    .Q(\data_array.data0[9][30] ));
 sky130_fd_sc_hd__dfxtp_2 _13606_ (.CLK(clk),
    .D(_02235_),
    .Q(\data_array.data0[9][31] ));
 sky130_fd_sc_hd__dfxtp_2 _13607_ (.CLK(clk),
    .D(_02236_),
    .Q(\data_array.data0[9][32] ));
 sky130_fd_sc_hd__dfxtp_2 _13608_ (.CLK(clk),
    .D(_02237_),
    .Q(\data_array.data0[9][33] ));
 sky130_fd_sc_hd__dfxtp_2 _13609_ (.CLK(clk),
    .D(_02238_),
    .Q(\data_array.data0[9][34] ));
 sky130_fd_sc_hd__dfxtp_2 _13610_ (.CLK(clk),
    .D(_02239_),
    .Q(\data_array.data0[9][35] ));
 sky130_fd_sc_hd__dfxtp_2 _13611_ (.CLK(clk),
    .D(_02240_),
    .Q(\data_array.data0[9][36] ));
 sky130_fd_sc_hd__dfxtp_2 _13612_ (.CLK(clk),
    .D(_02241_),
    .Q(\data_array.data0[9][37] ));
 sky130_fd_sc_hd__dfxtp_2 _13613_ (.CLK(clk),
    .D(_02242_),
    .Q(\data_array.data0[9][38] ));
 sky130_fd_sc_hd__dfxtp_2 _13614_ (.CLK(clk),
    .D(_02243_),
    .Q(\data_array.data0[9][39] ));
 sky130_fd_sc_hd__dfxtp_2 _13615_ (.CLK(clk),
    .D(_02244_),
    .Q(\data_array.data0[9][40] ));
 sky130_fd_sc_hd__dfxtp_2 _13616_ (.CLK(clk),
    .D(_02245_),
    .Q(\data_array.data0[9][41] ));
 sky130_fd_sc_hd__dfxtp_2 _13617_ (.CLK(clk),
    .D(_02246_),
    .Q(\data_array.data0[9][42] ));
 sky130_fd_sc_hd__dfxtp_2 _13618_ (.CLK(clk),
    .D(_02247_),
    .Q(\data_array.data0[9][43] ));
 sky130_fd_sc_hd__dfxtp_2 _13619_ (.CLK(clk),
    .D(_02248_),
    .Q(\data_array.data0[9][44] ));
 sky130_fd_sc_hd__dfxtp_2 _13620_ (.CLK(clk),
    .D(_02249_),
    .Q(\data_array.data0[9][45] ));
 sky130_fd_sc_hd__dfxtp_2 _13621_ (.CLK(clk),
    .D(_02250_),
    .Q(\data_array.data0[9][46] ));
 sky130_fd_sc_hd__dfxtp_2 _13622_ (.CLK(clk),
    .D(_02251_),
    .Q(\data_array.data0[9][47] ));
 sky130_fd_sc_hd__dfxtp_2 _13623_ (.CLK(clk),
    .D(_02252_),
    .Q(\data_array.data0[9][48] ));
 sky130_fd_sc_hd__dfxtp_2 _13624_ (.CLK(clk),
    .D(_02253_),
    .Q(\data_array.data0[9][49] ));
 sky130_fd_sc_hd__dfxtp_2 _13625_ (.CLK(clk),
    .D(_02254_),
    .Q(\data_array.data0[9][50] ));
 sky130_fd_sc_hd__dfxtp_2 _13626_ (.CLK(clk),
    .D(_02255_),
    .Q(\data_array.data0[9][51] ));
 sky130_fd_sc_hd__dfxtp_2 _13627_ (.CLK(clk),
    .D(_02256_),
    .Q(\data_array.data0[9][52] ));
 sky130_fd_sc_hd__dfxtp_2 _13628_ (.CLK(clk),
    .D(_02257_),
    .Q(\data_array.data0[9][53] ));
 sky130_fd_sc_hd__dfxtp_2 _13629_ (.CLK(clk),
    .D(_02258_),
    .Q(\data_array.data0[9][54] ));
 sky130_fd_sc_hd__dfxtp_2 _13630_ (.CLK(clk),
    .D(_02259_),
    .Q(\data_array.data0[9][55] ));
 sky130_fd_sc_hd__dfxtp_2 _13631_ (.CLK(clk),
    .D(_02260_),
    .Q(\data_array.data0[9][56] ));
 sky130_fd_sc_hd__dfxtp_2 _13632_ (.CLK(clk),
    .D(_02261_),
    .Q(\data_array.data0[9][57] ));
 sky130_fd_sc_hd__dfxtp_2 _13633_ (.CLK(clk),
    .D(_02262_),
    .Q(\data_array.data0[9][58] ));
 sky130_fd_sc_hd__dfxtp_2 _13634_ (.CLK(clk),
    .D(_02263_),
    .Q(\data_array.data0[9][59] ));
 sky130_fd_sc_hd__dfxtp_2 _13635_ (.CLK(clk),
    .D(_02264_),
    .Q(\data_array.data0[9][60] ));
 sky130_fd_sc_hd__dfxtp_2 _13636_ (.CLK(clk),
    .D(_02265_),
    .Q(\data_array.data0[9][61] ));
 sky130_fd_sc_hd__dfxtp_2 _13637_ (.CLK(clk),
    .D(_02266_),
    .Q(\data_array.data0[9][62] ));
 sky130_fd_sc_hd__dfxtp_2 _13638_ (.CLK(clk),
    .D(_02267_),
    .Q(\data_array.data0[9][63] ));
 sky130_fd_sc_hd__dfxtp_2 _13639_ (.CLK(clk),
    .D(_02268_),
    .Q(\tag_array.dirty0[9] ));
 sky130_fd_sc_hd__dfxtp_2 _13640_ (.CLK(clk),
    .D(_02269_),
    .Q(\data_array.data1[15][0] ));
 sky130_fd_sc_hd__dfxtp_2 _13641_ (.CLK(clk),
    .D(_02270_),
    .Q(\data_array.data1[15][1] ));
 sky130_fd_sc_hd__dfxtp_2 _13642_ (.CLK(clk),
    .D(_02271_),
    .Q(\data_array.data1[15][2] ));
 sky130_fd_sc_hd__dfxtp_2 _13643_ (.CLK(clk),
    .D(_02272_),
    .Q(\data_array.data1[15][3] ));
 sky130_fd_sc_hd__dfxtp_2 _13644_ (.CLK(clk),
    .D(_02273_),
    .Q(\data_array.data1[15][4] ));
 sky130_fd_sc_hd__dfxtp_2 _13645_ (.CLK(clk),
    .D(_02274_),
    .Q(\data_array.data1[15][5] ));
 sky130_fd_sc_hd__dfxtp_2 _13646_ (.CLK(clk),
    .D(_02275_),
    .Q(\data_array.data1[15][6] ));
 sky130_fd_sc_hd__dfxtp_2 _13647_ (.CLK(clk),
    .D(_02276_),
    .Q(\data_array.data1[15][7] ));
 sky130_fd_sc_hd__dfxtp_2 _13648_ (.CLK(clk),
    .D(_02277_),
    .Q(\data_array.data1[15][8] ));
 sky130_fd_sc_hd__dfxtp_2 _13649_ (.CLK(clk),
    .D(_02278_),
    .Q(\data_array.data1[15][9] ));
 sky130_fd_sc_hd__dfxtp_2 _13650_ (.CLK(clk),
    .D(_02279_),
    .Q(\data_array.data1[15][10] ));
 sky130_fd_sc_hd__dfxtp_2 _13651_ (.CLK(clk),
    .D(_02280_),
    .Q(\data_array.data1[15][11] ));
 sky130_fd_sc_hd__dfxtp_2 _13652_ (.CLK(clk),
    .D(_02281_),
    .Q(\data_array.data1[15][12] ));
 sky130_fd_sc_hd__dfxtp_2 _13653_ (.CLK(clk),
    .D(_02282_),
    .Q(\data_array.data1[15][13] ));
 sky130_fd_sc_hd__dfxtp_2 _13654_ (.CLK(clk),
    .D(_02283_),
    .Q(\data_array.data1[15][14] ));
 sky130_fd_sc_hd__dfxtp_2 _13655_ (.CLK(clk),
    .D(_02284_),
    .Q(\data_array.data1[15][15] ));
 sky130_fd_sc_hd__dfxtp_2 _13656_ (.CLK(clk),
    .D(_02285_),
    .Q(\data_array.data1[15][16] ));
 sky130_fd_sc_hd__dfxtp_2 _13657_ (.CLK(clk),
    .D(_02286_),
    .Q(\data_array.data1[15][17] ));
 sky130_fd_sc_hd__dfxtp_2 _13658_ (.CLK(clk),
    .D(_02287_),
    .Q(\data_array.data1[15][18] ));
 sky130_fd_sc_hd__dfxtp_2 _13659_ (.CLK(clk),
    .D(_02288_),
    .Q(\data_array.data1[15][19] ));
 sky130_fd_sc_hd__dfxtp_2 _13660_ (.CLK(clk),
    .D(_02289_),
    .Q(\data_array.data1[15][20] ));
 sky130_fd_sc_hd__dfxtp_2 _13661_ (.CLK(clk),
    .D(_02290_),
    .Q(\data_array.data1[15][21] ));
 sky130_fd_sc_hd__dfxtp_2 _13662_ (.CLK(clk),
    .D(_02291_),
    .Q(\data_array.data1[15][22] ));
 sky130_fd_sc_hd__dfxtp_2 _13663_ (.CLK(clk),
    .D(_02292_),
    .Q(\data_array.data1[15][23] ));
 sky130_fd_sc_hd__dfxtp_2 _13664_ (.CLK(clk),
    .D(_02293_),
    .Q(\data_array.data1[15][24] ));
 sky130_fd_sc_hd__dfxtp_2 _13665_ (.CLK(clk),
    .D(_02294_),
    .Q(\data_array.data1[15][25] ));
 sky130_fd_sc_hd__dfxtp_2 _13666_ (.CLK(clk),
    .D(_02295_),
    .Q(\data_array.data1[15][26] ));
 sky130_fd_sc_hd__dfxtp_2 _13667_ (.CLK(clk),
    .D(_02296_),
    .Q(\data_array.data1[15][27] ));
 sky130_fd_sc_hd__dfxtp_2 _13668_ (.CLK(clk),
    .D(_02297_),
    .Q(\data_array.data1[15][28] ));
 sky130_fd_sc_hd__dfxtp_2 _13669_ (.CLK(clk),
    .D(_02298_),
    .Q(\data_array.data1[15][29] ));
 sky130_fd_sc_hd__dfxtp_2 _13670_ (.CLK(clk),
    .D(_02299_),
    .Q(\data_array.data1[15][30] ));
 sky130_fd_sc_hd__dfxtp_2 _13671_ (.CLK(clk),
    .D(_02300_),
    .Q(\data_array.data1[15][31] ));
 sky130_fd_sc_hd__dfxtp_2 _13672_ (.CLK(clk),
    .D(_02301_),
    .Q(\data_array.data1[15][32] ));
 sky130_fd_sc_hd__dfxtp_2 _13673_ (.CLK(clk),
    .D(_02302_),
    .Q(\data_array.data1[15][33] ));
 sky130_fd_sc_hd__dfxtp_2 _13674_ (.CLK(clk),
    .D(_02303_),
    .Q(\data_array.data1[15][34] ));
 sky130_fd_sc_hd__dfxtp_2 _13675_ (.CLK(clk),
    .D(_02304_),
    .Q(\data_array.data1[15][35] ));
 sky130_fd_sc_hd__dfxtp_2 _13676_ (.CLK(clk),
    .D(_02305_),
    .Q(\data_array.data1[15][36] ));
 sky130_fd_sc_hd__dfxtp_2 _13677_ (.CLK(clk),
    .D(_02306_),
    .Q(\data_array.data1[15][37] ));
 sky130_fd_sc_hd__dfxtp_2 _13678_ (.CLK(clk),
    .D(_02307_),
    .Q(\data_array.data1[15][38] ));
 sky130_fd_sc_hd__dfxtp_2 _13679_ (.CLK(clk),
    .D(_02308_),
    .Q(\data_array.data1[15][39] ));
 sky130_fd_sc_hd__dfxtp_2 _13680_ (.CLK(clk),
    .D(_02309_),
    .Q(\data_array.data1[15][40] ));
 sky130_fd_sc_hd__dfxtp_2 _13681_ (.CLK(clk),
    .D(_02310_),
    .Q(\data_array.data1[15][41] ));
 sky130_fd_sc_hd__dfxtp_2 _13682_ (.CLK(clk),
    .D(_02311_),
    .Q(\data_array.data1[15][42] ));
 sky130_fd_sc_hd__dfxtp_2 _13683_ (.CLK(clk),
    .D(_02312_),
    .Q(\data_array.data1[15][43] ));
 sky130_fd_sc_hd__dfxtp_2 _13684_ (.CLK(clk),
    .D(_02313_),
    .Q(\data_array.data1[15][44] ));
 sky130_fd_sc_hd__dfxtp_2 _13685_ (.CLK(clk),
    .D(_02314_),
    .Q(\data_array.data1[15][45] ));
 sky130_fd_sc_hd__dfxtp_2 _13686_ (.CLK(clk),
    .D(_02315_),
    .Q(\data_array.data1[15][46] ));
 sky130_fd_sc_hd__dfxtp_2 _13687_ (.CLK(clk),
    .D(_02316_),
    .Q(\data_array.data1[15][47] ));
 sky130_fd_sc_hd__dfxtp_2 _13688_ (.CLK(clk),
    .D(_02317_),
    .Q(\data_array.data1[15][48] ));
 sky130_fd_sc_hd__dfxtp_2 _13689_ (.CLK(clk),
    .D(_02318_),
    .Q(\data_array.data1[15][49] ));
 sky130_fd_sc_hd__dfxtp_2 _13690_ (.CLK(clk),
    .D(_02319_),
    .Q(\data_array.data1[15][50] ));
 sky130_fd_sc_hd__dfxtp_2 _13691_ (.CLK(clk),
    .D(_02320_),
    .Q(\data_array.data1[15][51] ));
 sky130_fd_sc_hd__dfxtp_2 _13692_ (.CLK(clk),
    .D(_02321_),
    .Q(\data_array.data1[15][52] ));
 sky130_fd_sc_hd__dfxtp_2 _13693_ (.CLK(clk),
    .D(_02322_),
    .Q(\data_array.data1[15][53] ));
 sky130_fd_sc_hd__dfxtp_2 _13694_ (.CLK(clk),
    .D(_02323_),
    .Q(\data_array.data1[15][54] ));
 sky130_fd_sc_hd__dfxtp_2 _13695_ (.CLK(clk),
    .D(_02324_),
    .Q(\data_array.data1[15][55] ));
 sky130_fd_sc_hd__dfxtp_2 _13696_ (.CLK(clk),
    .D(_02325_),
    .Q(\data_array.data1[15][56] ));
 sky130_fd_sc_hd__dfxtp_2 _13697_ (.CLK(clk),
    .D(_02326_),
    .Q(\data_array.data1[15][57] ));
 sky130_fd_sc_hd__dfxtp_2 _13698_ (.CLK(clk),
    .D(_02327_),
    .Q(\data_array.data1[15][58] ));
 sky130_fd_sc_hd__dfxtp_2 _13699_ (.CLK(clk),
    .D(_02328_),
    .Q(\data_array.data1[15][59] ));
 sky130_fd_sc_hd__dfxtp_2 _13700_ (.CLK(clk),
    .D(_02329_),
    .Q(\data_array.data1[15][60] ));
 sky130_fd_sc_hd__dfxtp_2 _13701_ (.CLK(clk),
    .D(_02330_),
    .Q(\data_array.data1[15][61] ));
 sky130_fd_sc_hd__dfxtp_2 _13702_ (.CLK(clk),
    .D(_02331_),
    .Q(\data_array.data1[15][62] ));
 sky130_fd_sc_hd__dfxtp_2 _13703_ (.CLK(clk),
    .D(_02332_),
    .Q(\data_array.data1[15][63] ));
 sky130_fd_sc_hd__dfxtp_2 _13704_ (.CLK(clk),
    .D(_02333_),
    .Q(\data_array.data1[1][0] ));
 sky130_fd_sc_hd__dfxtp_2 _13705_ (.CLK(clk),
    .D(_02334_),
    .Q(\data_array.data1[1][1] ));
 sky130_fd_sc_hd__dfxtp_2 _13706_ (.CLK(clk),
    .D(_02335_),
    .Q(\data_array.data1[1][2] ));
 sky130_fd_sc_hd__dfxtp_2 _13707_ (.CLK(clk),
    .D(_02336_),
    .Q(\data_array.data1[1][3] ));
 sky130_fd_sc_hd__dfxtp_2 _13708_ (.CLK(clk),
    .D(_02337_),
    .Q(\data_array.data1[1][4] ));
 sky130_fd_sc_hd__dfxtp_2 _13709_ (.CLK(clk),
    .D(_02338_),
    .Q(\data_array.data1[1][5] ));
 sky130_fd_sc_hd__dfxtp_2 _13710_ (.CLK(clk),
    .D(_02339_),
    .Q(\data_array.data1[1][6] ));
 sky130_fd_sc_hd__dfxtp_2 _13711_ (.CLK(clk),
    .D(_02340_),
    .Q(\data_array.data1[1][7] ));
 sky130_fd_sc_hd__dfxtp_2 _13712_ (.CLK(clk),
    .D(_02341_),
    .Q(\data_array.data1[1][8] ));
 sky130_fd_sc_hd__dfxtp_2 _13713_ (.CLK(clk),
    .D(_02342_),
    .Q(\data_array.data1[1][9] ));
 sky130_fd_sc_hd__dfxtp_2 _13714_ (.CLK(clk),
    .D(_02343_),
    .Q(\data_array.data1[1][10] ));
 sky130_fd_sc_hd__dfxtp_2 _13715_ (.CLK(clk),
    .D(_02344_),
    .Q(\data_array.data1[1][11] ));
 sky130_fd_sc_hd__dfxtp_2 _13716_ (.CLK(clk),
    .D(_02345_),
    .Q(\data_array.data1[1][12] ));
 sky130_fd_sc_hd__dfxtp_2 _13717_ (.CLK(clk),
    .D(_02346_),
    .Q(\data_array.data1[1][13] ));
 sky130_fd_sc_hd__dfxtp_2 _13718_ (.CLK(clk),
    .D(_02347_),
    .Q(\data_array.data1[1][14] ));
 sky130_fd_sc_hd__dfxtp_2 _13719_ (.CLK(clk),
    .D(_02348_),
    .Q(\data_array.data1[1][15] ));
 sky130_fd_sc_hd__dfxtp_2 _13720_ (.CLK(clk),
    .D(_02349_),
    .Q(\data_array.data1[1][16] ));
 sky130_fd_sc_hd__dfxtp_2 _13721_ (.CLK(clk),
    .D(_02350_),
    .Q(\data_array.data1[1][17] ));
 sky130_fd_sc_hd__dfxtp_2 _13722_ (.CLK(clk),
    .D(_02351_),
    .Q(\data_array.data1[1][18] ));
 sky130_fd_sc_hd__dfxtp_2 _13723_ (.CLK(clk),
    .D(_02352_),
    .Q(\data_array.data1[1][19] ));
 sky130_fd_sc_hd__dfxtp_2 _13724_ (.CLK(clk),
    .D(_02353_),
    .Q(\data_array.data1[1][20] ));
 sky130_fd_sc_hd__dfxtp_2 _13725_ (.CLK(clk),
    .D(_02354_),
    .Q(\data_array.data1[1][21] ));
 sky130_fd_sc_hd__dfxtp_2 _13726_ (.CLK(clk),
    .D(_02355_),
    .Q(\data_array.data1[1][22] ));
 sky130_fd_sc_hd__dfxtp_2 _13727_ (.CLK(clk),
    .D(_02356_),
    .Q(\data_array.data1[1][23] ));
 sky130_fd_sc_hd__dfxtp_2 _13728_ (.CLK(clk),
    .D(_02357_),
    .Q(\data_array.data1[1][24] ));
 sky130_fd_sc_hd__dfxtp_2 _13729_ (.CLK(clk),
    .D(_02358_),
    .Q(\data_array.data1[1][25] ));
 sky130_fd_sc_hd__dfxtp_2 _13730_ (.CLK(clk),
    .D(_02359_),
    .Q(\data_array.data1[1][26] ));
 sky130_fd_sc_hd__dfxtp_2 _13731_ (.CLK(clk),
    .D(_02360_),
    .Q(\data_array.data1[1][27] ));
 sky130_fd_sc_hd__dfxtp_2 _13732_ (.CLK(clk),
    .D(_02361_),
    .Q(\data_array.data1[1][28] ));
 sky130_fd_sc_hd__dfxtp_2 _13733_ (.CLK(clk),
    .D(_02362_),
    .Q(\data_array.data1[1][29] ));
 sky130_fd_sc_hd__dfxtp_2 _13734_ (.CLK(clk),
    .D(_02363_),
    .Q(\data_array.data1[1][30] ));
 sky130_fd_sc_hd__dfxtp_2 _13735_ (.CLK(clk),
    .D(_02364_),
    .Q(\data_array.data1[1][31] ));
 sky130_fd_sc_hd__dfxtp_2 _13736_ (.CLK(clk),
    .D(_02365_),
    .Q(\data_array.data1[1][32] ));
 sky130_fd_sc_hd__dfxtp_2 _13737_ (.CLK(clk),
    .D(_02366_),
    .Q(\data_array.data1[1][33] ));
 sky130_fd_sc_hd__dfxtp_2 _13738_ (.CLK(clk),
    .D(_02367_),
    .Q(\data_array.data1[1][34] ));
 sky130_fd_sc_hd__dfxtp_2 _13739_ (.CLK(clk),
    .D(_02368_),
    .Q(\data_array.data1[1][35] ));
 sky130_fd_sc_hd__dfxtp_2 _13740_ (.CLK(clk),
    .D(_02369_),
    .Q(\data_array.data1[1][36] ));
 sky130_fd_sc_hd__dfxtp_2 _13741_ (.CLK(clk),
    .D(_02370_),
    .Q(\data_array.data1[1][37] ));
 sky130_fd_sc_hd__dfxtp_2 _13742_ (.CLK(clk),
    .D(_02371_),
    .Q(\data_array.data1[1][38] ));
 sky130_fd_sc_hd__dfxtp_2 _13743_ (.CLK(clk),
    .D(_02372_),
    .Q(\data_array.data1[1][39] ));
 sky130_fd_sc_hd__dfxtp_2 _13744_ (.CLK(clk),
    .D(_02373_),
    .Q(\data_array.data1[1][40] ));
 sky130_fd_sc_hd__dfxtp_2 _13745_ (.CLK(clk),
    .D(_02374_),
    .Q(\data_array.data1[1][41] ));
 sky130_fd_sc_hd__dfxtp_2 _13746_ (.CLK(clk),
    .D(_02375_),
    .Q(\data_array.data1[1][42] ));
 sky130_fd_sc_hd__dfxtp_2 _13747_ (.CLK(clk),
    .D(_02376_),
    .Q(\data_array.data1[1][43] ));
 sky130_fd_sc_hd__dfxtp_2 _13748_ (.CLK(clk),
    .D(_02377_),
    .Q(\data_array.data1[1][44] ));
 sky130_fd_sc_hd__dfxtp_2 _13749_ (.CLK(clk),
    .D(_02378_),
    .Q(\data_array.data1[1][45] ));
 sky130_fd_sc_hd__dfxtp_2 _13750_ (.CLK(clk),
    .D(_02379_),
    .Q(\data_array.data1[1][46] ));
 sky130_fd_sc_hd__dfxtp_2 _13751_ (.CLK(clk),
    .D(_02380_),
    .Q(\data_array.data1[1][47] ));
 sky130_fd_sc_hd__dfxtp_2 _13752_ (.CLK(clk),
    .D(_02381_),
    .Q(\data_array.data1[1][48] ));
 sky130_fd_sc_hd__dfxtp_2 _13753_ (.CLK(clk),
    .D(_02382_),
    .Q(\data_array.data1[1][49] ));
 sky130_fd_sc_hd__dfxtp_2 _13754_ (.CLK(clk),
    .D(_02383_),
    .Q(\data_array.data1[1][50] ));
 sky130_fd_sc_hd__dfxtp_2 _13755_ (.CLK(clk),
    .D(_02384_),
    .Q(\data_array.data1[1][51] ));
 sky130_fd_sc_hd__dfxtp_2 _13756_ (.CLK(clk),
    .D(_02385_),
    .Q(\data_array.data1[1][52] ));
 sky130_fd_sc_hd__dfxtp_2 _13757_ (.CLK(clk),
    .D(_02386_),
    .Q(\data_array.data1[1][53] ));
 sky130_fd_sc_hd__dfxtp_2 _13758_ (.CLK(clk),
    .D(_02387_),
    .Q(\data_array.data1[1][54] ));
 sky130_fd_sc_hd__dfxtp_2 _13759_ (.CLK(clk),
    .D(_02388_),
    .Q(\data_array.data1[1][55] ));
 sky130_fd_sc_hd__dfxtp_2 _13760_ (.CLK(clk),
    .D(_02389_),
    .Q(\data_array.data1[1][56] ));
 sky130_fd_sc_hd__dfxtp_2 _13761_ (.CLK(clk),
    .D(_02390_),
    .Q(\data_array.data1[1][57] ));
 sky130_fd_sc_hd__dfxtp_2 _13762_ (.CLK(clk),
    .D(_02391_),
    .Q(\data_array.data1[1][58] ));
 sky130_fd_sc_hd__dfxtp_2 _13763_ (.CLK(clk),
    .D(_02392_),
    .Q(\data_array.data1[1][59] ));
 sky130_fd_sc_hd__dfxtp_2 _13764_ (.CLK(clk),
    .D(_02393_),
    .Q(\data_array.data1[1][60] ));
 sky130_fd_sc_hd__dfxtp_2 _13765_ (.CLK(clk),
    .D(_02394_),
    .Q(\data_array.data1[1][61] ));
 sky130_fd_sc_hd__dfxtp_2 _13766_ (.CLK(clk),
    .D(_02395_),
    .Q(\data_array.data1[1][62] ));
 sky130_fd_sc_hd__dfxtp_2 _13767_ (.CLK(clk),
    .D(_02396_),
    .Q(\data_array.data1[1][63] ));
 sky130_fd_sc_hd__dfxtp_2 _13768_ (.CLK(clk),
    .D(_02397_),
    .Q(\data_array.data1[2][0] ));
 sky130_fd_sc_hd__dfxtp_2 _13769_ (.CLK(clk),
    .D(_02398_),
    .Q(\data_array.data1[2][1] ));
 sky130_fd_sc_hd__dfxtp_2 _13770_ (.CLK(clk),
    .D(_02399_),
    .Q(\data_array.data1[2][2] ));
 sky130_fd_sc_hd__dfxtp_2 _13771_ (.CLK(clk),
    .D(_02400_),
    .Q(\data_array.data1[2][3] ));
 sky130_fd_sc_hd__dfxtp_2 _13772_ (.CLK(clk),
    .D(_02401_),
    .Q(\data_array.data1[2][4] ));
 sky130_fd_sc_hd__dfxtp_2 _13773_ (.CLK(clk),
    .D(_02402_),
    .Q(\data_array.data1[2][5] ));
 sky130_fd_sc_hd__dfxtp_2 _13774_ (.CLK(clk),
    .D(_02403_),
    .Q(\data_array.data1[2][6] ));
 sky130_fd_sc_hd__dfxtp_2 _13775_ (.CLK(clk),
    .D(_02404_),
    .Q(\data_array.data1[2][7] ));
 sky130_fd_sc_hd__dfxtp_2 _13776_ (.CLK(clk),
    .D(_02405_),
    .Q(\data_array.data1[2][8] ));
 sky130_fd_sc_hd__dfxtp_2 _13777_ (.CLK(clk),
    .D(_02406_),
    .Q(\data_array.data1[2][9] ));
 sky130_fd_sc_hd__dfxtp_2 _13778_ (.CLK(clk),
    .D(_02407_),
    .Q(\data_array.data1[2][10] ));
 sky130_fd_sc_hd__dfxtp_2 _13779_ (.CLK(clk),
    .D(_02408_),
    .Q(\data_array.data1[2][11] ));
 sky130_fd_sc_hd__dfxtp_2 _13780_ (.CLK(clk),
    .D(_02409_),
    .Q(\data_array.data1[2][12] ));
 sky130_fd_sc_hd__dfxtp_2 _13781_ (.CLK(clk),
    .D(_02410_),
    .Q(\data_array.data1[2][13] ));
 sky130_fd_sc_hd__dfxtp_2 _13782_ (.CLK(clk),
    .D(_02411_),
    .Q(\data_array.data1[2][14] ));
 sky130_fd_sc_hd__dfxtp_2 _13783_ (.CLK(clk),
    .D(_02412_),
    .Q(\data_array.data1[2][15] ));
 sky130_fd_sc_hd__dfxtp_2 _13784_ (.CLK(clk),
    .D(_02413_),
    .Q(\data_array.data1[2][16] ));
 sky130_fd_sc_hd__dfxtp_2 _13785_ (.CLK(clk),
    .D(_02414_),
    .Q(\data_array.data1[2][17] ));
 sky130_fd_sc_hd__dfxtp_2 _13786_ (.CLK(clk),
    .D(_02415_),
    .Q(\data_array.data1[2][18] ));
 sky130_fd_sc_hd__dfxtp_2 _13787_ (.CLK(clk),
    .D(_02416_),
    .Q(\data_array.data1[2][19] ));
 sky130_fd_sc_hd__dfxtp_2 _13788_ (.CLK(clk),
    .D(_02417_),
    .Q(\data_array.data1[2][20] ));
 sky130_fd_sc_hd__dfxtp_2 _13789_ (.CLK(clk),
    .D(_02418_),
    .Q(\data_array.data1[2][21] ));
 sky130_fd_sc_hd__dfxtp_2 _13790_ (.CLK(clk),
    .D(_02419_),
    .Q(\data_array.data1[2][22] ));
 sky130_fd_sc_hd__dfxtp_2 _13791_ (.CLK(clk),
    .D(_02420_),
    .Q(\data_array.data1[2][23] ));
 sky130_fd_sc_hd__dfxtp_2 _13792_ (.CLK(clk),
    .D(_02421_),
    .Q(\data_array.data1[2][24] ));
 sky130_fd_sc_hd__dfxtp_2 _13793_ (.CLK(clk),
    .D(_02422_),
    .Q(\data_array.data1[2][25] ));
 sky130_fd_sc_hd__dfxtp_2 _13794_ (.CLK(clk),
    .D(_02423_),
    .Q(\data_array.data1[2][26] ));
 sky130_fd_sc_hd__dfxtp_2 _13795_ (.CLK(clk),
    .D(_02424_),
    .Q(\data_array.data1[2][27] ));
 sky130_fd_sc_hd__dfxtp_2 _13796_ (.CLK(clk),
    .D(_02425_),
    .Q(\data_array.data1[2][28] ));
 sky130_fd_sc_hd__dfxtp_2 _13797_ (.CLK(clk),
    .D(_02426_),
    .Q(\data_array.data1[2][29] ));
 sky130_fd_sc_hd__dfxtp_2 _13798_ (.CLK(clk),
    .D(_02427_),
    .Q(\data_array.data1[2][30] ));
 sky130_fd_sc_hd__dfxtp_2 _13799_ (.CLK(clk),
    .D(_02428_),
    .Q(\data_array.data1[2][31] ));
 sky130_fd_sc_hd__dfxtp_2 _13800_ (.CLK(clk),
    .D(_02429_),
    .Q(\data_array.data1[2][32] ));
 sky130_fd_sc_hd__dfxtp_2 _13801_ (.CLK(clk),
    .D(_02430_),
    .Q(\data_array.data1[2][33] ));
 sky130_fd_sc_hd__dfxtp_2 _13802_ (.CLK(clk),
    .D(_02431_),
    .Q(\data_array.data1[2][34] ));
 sky130_fd_sc_hd__dfxtp_2 _13803_ (.CLK(clk),
    .D(_02432_),
    .Q(\data_array.data1[2][35] ));
 sky130_fd_sc_hd__dfxtp_2 _13804_ (.CLK(clk),
    .D(_02433_),
    .Q(\data_array.data1[2][36] ));
 sky130_fd_sc_hd__dfxtp_2 _13805_ (.CLK(clk),
    .D(_02434_),
    .Q(\data_array.data1[2][37] ));
 sky130_fd_sc_hd__dfxtp_2 _13806_ (.CLK(clk),
    .D(_02435_),
    .Q(\data_array.data1[2][38] ));
 sky130_fd_sc_hd__dfxtp_2 _13807_ (.CLK(clk),
    .D(_02436_),
    .Q(\data_array.data1[2][39] ));
 sky130_fd_sc_hd__dfxtp_2 _13808_ (.CLK(clk),
    .D(_02437_),
    .Q(\data_array.data1[2][40] ));
 sky130_fd_sc_hd__dfxtp_2 _13809_ (.CLK(clk),
    .D(_02438_),
    .Q(\data_array.data1[2][41] ));
 sky130_fd_sc_hd__dfxtp_2 _13810_ (.CLK(clk),
    .D(_02439_),
    .Q(\data_array.data1[2][42] ));
 sky130_fd_sc_hd__dfxtp_2 _13811_ (.CLK(clk),
    .D(_02440_),
    .Q(\data_array.data1[2][43] ));
 sky130_fd_sc_hd__dfxtp_2 _13812_ (.CLK(clk),
    .D(_02441_),
    .Q(\data_array.data1[2][44] ));
 sky130_fd_sc_hd__dfxtp_2 _13813_ (.CLK(clk),
    .D(_02442_),
    .Q(\data_array.data1[2][45] ));
 sky130_fd_sc_hd__dfxtp_2 _13814_ (.CLK(clk),
    .D(_02443_),
    .Q(\data_array.data1[2][46] ));
 sky130_fd_sc_hd__dfxtp_2 _13815_ (.CLK(clk),
    .D(_02444_),
    .Q(\data_array.data1[2][47] ));
 sky130_fd_sc_hd__dfxtp_2 _13816_ (.CLK(clk),
    .D(_02445_),
    .Q(\data_array.data1[2][48] ));
 sky130_fd_sc_hd__dfxtp_2 _13817_ (.CLK(clk),
    .D(_02446_),
    .Q(\data_array.data1[2][49] ));
 sky130_fd_sc_hd__dfxtp_2 _13818_ (.CLK(clk),
    .D(_02447_),
    .Q(\data_array.data1[2][50] ));
 sky130_fd_sc_hd__dfxtp_2 _13819_ (.CLK(clk),
    .D(_02448_),
    .Q(\data_array.data1[2][51] ));
 sky130_fd_sc_hd__dfxtp_2 _13820_ (.CLK(clk),
    .D(_02449_),
    .Q(\data_array.data1[2][52] ));
 sky130_fd_sc_hd__dfxtp_2 _13821_ (.CLK(clk),
    .D(_02450_),
    .Q(\data_array.data1[2][53] ));
 sky130_fd_sc_hd__dfxtp_2 _13822_ (.CLK(clk),
    .D(_02451_),
    .Q(\data_array.data1[2][54] ));
 sky130_fd_sc_hd__dfxtp_2 _13823_ (.CLK(clk),
    .D(_02452_),
    .Q(\data_array.data1[2][55] ));
 sky130_fd_sc_hd__dfxtp_2 _13824_ (.CLK(clk),
    .D(_02453_),
    .Q(\data_array.data1[2][56] ));
 sky130_fd_sc_hd__dfxtp_2 _13825_ (.CLK(clk),
    .D(_02454_),
    .Q(\data_array.data1[2][57] ));
 sky130_fd_sc_hd__dfxtp_2 _13826_ (.CLK(clk),
    .D(_02455_),
    .Q(\data_array.data1[2][58] ));
 sky130_fd_sc_hd__dfxtp_2 _13827_ (.CLK(clk),
    .D(_02456_),
    .Q(\data_array.data1[2][59] ));
 sky130_fd_sc_hd__dfxtp_2 _13828_ (.CLK(clk),
    .D(_02457_),
    .Q(\data_array.data1[2][60] ));
 sky130_fd_sc_hd__dfxtp_2 _13829_ (.CLK(clk),
    .D(_02458_),
    .Q(\data_array.data1[2][61] ));
 sky130_fd_sc_hd__dfxtp_2 _13830_ (.CLK(clk),
    .D(_02459_),
    .Q(\data_array.data1[2][62] ));
 sky130_fd_sc_hd__dfxtp_2 _13831_ (.CLK(clk),
    .D(_02460_),
    .Q(\data_array.data1[2][63] ));
 sky130_fd_sc_hd__dfxtp_2 _13832_ (.CLK(clk),
    .D(_02461_),
    .Q(\data_array.data1[3][0] ));
 sky130_fd_sc_hd__dfxtp_2 _13833_ (.CLK(clk),
    .D(_02462_),
    .Q(\data_array.data1[3][1] ));
 sky130_fd_sc_hd__dfxtp_2 _13834_ (.CLK(clk),
    .D(_02463_),
    .Q(\data_array.data1[3][2] ));
 sky130_fd_sc_hd__dfxtp_2 _13835_ (.CLK(clk),
    .D(_02464_),
    .Q(\data_array.data1[3][3] ));
 sky130_fd_sc_hd__dfxtp_2 _13836_ (.CLK(clk),
    .D(_02465_),
    .Q(\data_array.data1[3][4] ));
 sky130_fd_sc_hd__dfxtp_2 _13837_ (.CLK(clk),
    .D(_02466_),
    .Q(\data_array.data1[3][5] ));
 sky130_fd_sc_hd__dfxtp_2 _13838_ (.CLK(clk),
    .D(_02467_),
    .Q(\data_array.data1[3][6] ));
 sky130_fd_sc_hd__dfxtp_2 _13839_ (.CLK(clk),
    .D(_02468_),
    .Q(\data_array.data1[3][7] ));
 sky130_fd_sc_hd__dfxtp_2 _13840_ (.CLK(clk),
    .D(_02469_),
    .Q(\data_array.data1[3][8] ));
 sky130_fd_sc_hd__dfxtp_2 _13841_ (.CLK(clk),
    .D(_02470_),
    .Q(\data_array.data1[3][9] ));
 sky130_fd_sc_hd__dfxtp_2 _13842_ (.CLK(clk),
    .D(_02471_),
    .Q(\data_array.data1[3][10] ));
 sky130_fd_sc_hd__dfxtp_2 _13843_ (.CLK(clk),
    .D(_02472_),
    .Q(\data_array.data1[3][11] ));
 sky130_fd_sc_hd__dfxtp_2 _13844_ (.CLK(clk),
    .D(_02473_),
    .Q(\data_array.data1[3][12] ));
 sky130_fd_sc_hd__dfxtp_2 _13845_ (.CLK(clk),
    .D(_02474_),
    .Q(\data_array.data1[3][13] ));
 sky130_fd_sc_hd__dfxtp_2 _13846_ (.CLK(clk),
    .D(_02475_),
    .Q(\data_array.data1[3][14] ));
 sky130_fd_sc_hd__dfxtp_2 _13847_ (.CLK(clk),
    .D(_02476_),
    .Q(\data_array.data1[3][15] ));
 sky130_fd_sc_hd__dfxtp_2 _13848_ (.CLK(clk),
    .D(_02477_),
    .Q(\data_array.data1[3][16] ));
 sky130_fd_sc_hd__dfxtp_2 _13849_ (.CLK(clk),
    .D(_02478_),
    .Q(\data_array.data1[3][17] ));
 sky130_fd_sc_hd__dfxtp_2 _13850_ (.CLK(clk),
    .D(_02479_),
    .Q(\data_array.data1[3][18] ));
 sky130_fd_sc_hd__dfxtp_2 _13851_ (.CLK(clk),
    .D(_02480_),
    .Q(\data_array.data1[3][19] ));
 sky130_fd_sc_hd__dfxtp_2 _13852_ (.CLK(clk),
    .D(_02481_),
    .Q(\data_array.data1[3][20] ));
 sky130_fd_sc_hd__dfxtp_2 _13853_ (.CLK(clk),
    .D(_02482_),
    .Q(\data_array.data1[3][21] ));
 sky130_fd_sc_hd__dfxtp_2 _13854_ (.CLK(clk),
    .D(_02483_),
    .Q(\data_array.data1[3][22] ));
 sky130_fd_sc_hd__dfxtp_2 _13855_ (.CLK(clk),
    .D(_02484_),
    .Q(\data_array.data1[3][23] ));
 sky130_fd_sc_hd__dfxtp_2 _13856_ (.CLK(clk),
    .D(_02485_),
    .Q(\data_array.data1[3][24] ));
 sky130_fd_sc_hd__dfxtp_2 _13857_ (.CLK(clk),
    .D(_02486_),
    .Q(\data_array.data1[3][25] ));
 sky130_fd_sc_hd__dfxtp_2 _13858_ (.CLK(clk),
    .D(_02487_),
    .Q(\data_array.data1[3][26] ));
 sky130_fd_sc_hd__dfxtp_2 _13859_ (.CLK(clk),
    .D(_02488_),
    .Q(\data_array.data1[3][27] ));
 sky130_fd_sc_hd__dfxtp_2 _13860_ (.CLK(clk),
    .D(_02489_),
    .Q(\data_array.data1[3][28] ));
 sky130_fd_sc_hd__dfxtp_2 _13861_ (.CLK(clk),
    .D(_02490_),
    .Q(\data_array.data1[3][29] ));
 sky130_fd_sc_hd__dfxtp_2 _13862_ (.CLK(clk),
    .D(_02491_),
    .Q(\data_array.data1[3][30] ));
 sky130_fd_sc_hd__dfxtp_2 _13863_ (.CLK(clk),
    .D(_02492_),
    .Q(\data_array.data1[3][31] ));
 sky130_fd_sc_hd__dfxtp_2 _13864_ (.CLK(clk),
    .D(_02493_),
    .Q(\data_array.data1[3][32] ));
 sky130_fd_sc_hd__dfxtp_2 _13865_ (.CLK(clk),
    .D(_02494_),
    .Q(\data_array.data1[3][33] ));
 sky130_fd_sc_hd__dfxtp_2 _13866_ (.CLK(clk),
    .D(_02495_),
    .Q(\data_array.data1[3][34] ));
 sky130_fd_sc_hd__dfxtp_2 _13867_ (.CLK(clk),
    .D(_02496_),
    .Q(\data_array.data1[3][35] ));
 sky130_fd_sc_hd__dfxtp_2 _13868_ (.CLK(clk),
    .D(_02497_),
    .Q(\data_array.data1[3][36] ));
 sky130_fd_sc_hd__dfxtp_2 _13869_ (.CLK(clk),
    .D(_02498_),
    .Q(\data_array.data1[3][37] ));
 sky130_fd_sc_hd__dfxtp_2 _13870_ (.CLK(clk),
    .D(_02499_),
    .Q(\data_array.data1[3][38] ));
 sky130_fd_sc_hd__dfxtp_2 _13871_ (.CLK(clk),
    .D(_02500_),
    .Q(\data_array.data1[3][39] ));
 sky130_fd_sc_hd__dfxtp_2 _13872_ (.CLK(clk),
    .D(_02501_),
    .Q(\data_array.data1[3][40] ));
 sky130_fd_sc_hd__dfxtp_2 _13873_ (.CLK(clk),
    .D(_02502_),
    .Q(\data_array.data1[3][41] ));
 sky130_fd_sc_hd__dfxtp_2 _13874_ (.CLK(clk),
    .D(_02503_),
    .Q(\data_array.data1[3][42] ));
 sky130_fd_sc_hd__dfxtp_2 _13875_ (.CLK(clk),
    .D(_02504_),
    .Q(\data_array.data1[3][43] ));
 sky130_fd_sc_hd__dfxtp_2 _13876_ (.CLK(clk),
    .D(_02505_),
    .Q(\data_array.data1[3][44] ));
 sky130_fd_sc_hd__dfxtp_2 _13877_ (.CLK(clk),
    .D(_02506_),
    .Q(\data_array.data1[3][45] ));
 sky130_fd_sc_hd__dfxtp_2 _13878_ (.CLK(clk),
    .D(_02507_),
    .Q(\data_array.data1[3][46] ));
 sky130_fd_sc_hd__dfxtp_2 _13879_ (.CLK(clk),
    .D(_02508_),
    .Q(\data_array.data1[3][47] ));
 sky130_fd_sc_hd__dfxtp_2 _13880_ (.CLK(clk),
    .D(_02509_),
    .Q(\data_array.data1[3][48] ));
 sky130_fd_sc_hd__dfxtp_2 _13881_ (.CLK(clk),
    .D(_02510_),
    .Q(\data_array.data1[3][49] ));
 sky130_fd_sc_hd__dfxtp_2 _13882_ (.CLK(clk),
    .D(_02511_),
    .Q(\data_array.data1[3][50] ));
 sky130_fd_sc_hd__dfxtp_2 _13883_ (.CLK(clk),
    .D(_02512_),
    .Q(\data_array.data1[3][51] ));
 sky130_fd_sc_hd__dfxtp_2 _13884_ (.CLK(clk),
    .D(_02513_),
    .Q(\data_array.data1[3][52] ));
 sky130_fd_sc_hd__dfxtp_2 _13885_ (.CLK(clk),
    .D(_02514_),
    .Q(\data_array.data1[3][53] ));
 sky130_fd_sc_hd__dfxtp_2 _13886_ (.CLK(clk),
    .D(_02515_),
    .Q(\data_array.data1[3][54] ));
 sky130_fd_sc_hd__dfxtp_2 _13887_ (.CLK(clk),
    .D(_02516_),
    .Q(\data_array.data1[3][55] ));
 sky130_fd_sc_hd__dfxtp_2 _13888_ (.CLK(clk),
    .D(_02517_),
    .Q(\data_array.data1[3][56] ));
 sky130_fd_sc_hd__dfxtp_2 _13889_ (.CLK(clk),
    .D(_02518_),
    .Q(\data_array.data1[3][57] ));
 sky130_fd_sc_hd__dfxtp_2 _13890_ (.CLK(clk),
    .D(_02519_),
    .Q(\data_array.data1[3][58] ));
 sky130_fd_sc_hd__dfxtp_2 _13891_ (.CLK(clk),
    .D(_02520_),
    .Q(\data_array.data1[3][59] ));
 sky130_fd_sc_hd__dfxtp_2 _13892_ (.CLK(clk),
    .D(_02521_),
    .Q(\data_array.data1[3][60] ));
 sky130_fd_sc_hd__dfxtp_2 _13893_ (.CLK(clk),
    .D(_02522_),
    .Q(\data_array.data1[3][61] ));
 sky130_fd_sc_hd__dfxtp_2 _13894_ (.CLK(clk),
    .D(_02523_),
    .Q(\data_array.data1[3][62] ));
 sky130_fd_sc_hd__dfxtp_2 _13895_ (.CLK(clk),
    .D(_02524_),
    .Q(\data_array.data1[3][63] ));
 sky130_fd_sc_hd__dfxtp_2 _13896_ (.CLK(clk),
    .D(_02525_),
    .Q(\data_array.data1[4][0] ));
 sky130_fd_sc_hd__dfxtp_2 _13897_ (.CLK(clk),
    .D(_02526_),
    .Q(\data_array.data1[4][1] ));
 sky130_fd_sc_hd__dfxtp_2 _13898_ (.CLK(clk),
    .D(_02527_),
    .Q(\data_array.data1[4][2] ));
 sky130_fd_sc_hd__dfxtp_2 _13899_ (.CLK(clk),
    .D(_02528_),
    .Q(\data_array.data1[4][3] ));
 sky130_fd_sc_hd__dfxtp_2 _13900_ (.CLK(clk),
    .D(_02529_),
    .Q(\data_array.data1[4][4] ));
 sky130_fd_sc_hd__dfxtp_2 _13901_ (.CLK(clk),
    .D(_02530_),
    .Q(\data_array.data1[4][5] ));
 sky130_fd_sc_hd__dfxtp_2 _13902_ (.CLK(clk),
    .D(_02531_),
    .Q(\data_array.data1[4][6] ));
 sky130_fd_sc_hd__dfxtp_2 _13903_ (.CLK(clk),
    .D(_02532_),
    .Q(\data_array.data1[4][7] ));
 sky130_fd_sc_hd__dfxtp_2 _13904_ (.CLK(clk),
    .D(_02533_),
    .Q(\data_array.data1[4][8] ));
 sky130_fd_sc_hd__dfxtp_2 _13905_ (.CLK(clk),
    .D(_02534_),
    .Q(\data_array.data1[4][9] ));
 sky130_fd_sc_hd__dfxtp_2 _13906_ (.CLK(clk),
    .D(_02535_),
    .Q(\data_array.data1[4][10] ));
 sky130_fd_sc_hd__dfxtp_2 _13907_ (.CLK(clk),
    .D(_02536_),
    .Q(\data_array.data1[4][11] ));
 sky130_fd_sc_hd__dfxtp_2 _13908_ (.CLK(clk),
    .D(_02537_),
    .Q(\data_array.data1[4][12] ));
 sky130_fd_sc_hd__dfxtp_2 _13909_ (.CLK(clk),
    .D(_02538_),
    .Q(\data_array.data1[4][13] ));
 sky130_fd_sc_hd__dfxtp_2 _13910_ (.CLK(clk),
    .D(_02539_),
    .Q(\data_array.data1[4][14] ));
 sky130_fd_sc_hd__dfxtp_2 _13911_ (.CLK(clk),
    .D(_02540_),
    .Q(\data_array.data1[4][15] ));
 sky130_fd_sc_hd__dfxtp_2 _13912_ (.CLK(clk),
    .D(_02541_),
    .Q(\data_array.data1[4][16] ));
 sky130_fd_sc_hd__dfxtp_2 _13913_ (.CLK(clk),
    .D(_02542_),
    .Q(\data_array.data1[4][17] ));
 sky130_fd_sc_hd__dfxtp_2 _13914_ (.CLK(clk),
    .D(_02543_),
    .Q(\data_array.data1[4][18] ));
 sky130_fd_sc_hd__dfxtp_2 _13915_ (.CLK(clk),
    .D(_02544_),
    .Q(\data_array.data1[4][19] ));
 sky130_fd_sc_hd__dfxtp_2 _13916_ (.CLK(clk),
    .D(_02545_),
    .Q(\data_array.data1[4][20] ));
 sky130_fd_sc_hd__dfxtp_2 _13917_ (.CLK(clk),
    .D(_02546_),
    .Q(\data_array.data1[4][21] ));
 sky130_fd_sc_hd__dfxtp_2 _13918_ (.CLK(clk),
    .D(_02547_),
    .Q(\data_array.data1[4][22] ));
 sky130_fd_sc_hd__dfxtp_2 _13919_ (.CLK(clk),
    .D(_02548_),
    .Q(\data_array.data1[4][23] ));
 sky130_fd_sc_hd__dfxtp_2 _13920_ (.CLK(clk),
    .D(_02549_),
    .Q(\data_array.data1[4][24] ));
 sky130_fd_sc_hd__dfxtp_2 _13921_ (.CLK(clk),
    .D(_02550_),
    .Q(\data_array.data1[4][25] ));
 sky130_fd_sc_hd__dfxtp_2 _13922_ (.CLK(clk),
    .D(_02551_),
    .Q(\data_array.data1[4][26] ));
 sky130_fd_sc_hd__dfxtp_2 _13923_ (.CLK(clk),
    .D(_02552_),
    .Q(\data_array.data1[4][27] ));
 sky130_fd_sc_hd__dfxtp_2 _13924_ (.CLK(clk),
    .D(_02553_),
    .Q(\data_array.data1[4][28] ));
 sky130_fd_sc_hd__dfxtp_2 _13925_ (.CLK(clk),
    .D(_02554_),
    .Q(\data_array.data1[4][29] ));
 sky130_fd_sc_hd__dfxtp_2 _13926_ (.CLK(clk),
    .D(_02555_),
    .Q(\data_array.data1[4][30] ));
 sky130_fd_sc_hd__dfxtp_2 _13927_ (.CLK(clk),
    .D(_02556_),
    .Q(\data_array.data1[4][31] ));
 sky130_fd_sc_hd__dfxtp_2 _13928_ (.CLK(clk),
    .D(_02557_),
    .Q(\data_array.data1[4][32] ));
 sky130_fd_sc_hd__dfxtp_2 _13929_ (.CLK(clk),
    .D(_02558_),
    .Q(\data_array.data1[4][33] ));
 sky130_fd_sc_hd__dfxtp_2 _13930_ (.CLK(clk),
    .D(_02559_),
    .Q(\data_array.data1[4][34] ));
 sky130_fd_sc_hd__dfxtp_2 _13931_ (.CLK(clk),
    .D(_02560_),
    .Q(\data_array.data1[4][35] ));
 sky130_fd_sc_hd__dfxtp_2 _13932_ (.CLK(clk),
    .D(_02561_),
    .Q(\data_array.data1[4][36] ));
 sky130_fd_sc_hd__dfxtp_2 _13933_ (.CLK(clk),
    .D(_02562_),
    .Q(\data_array.data1[4][37] ));
 sky130_fd_sc_hd__dfxtp_2 _13934_ (.CLK(clk),
    .D(_02563_),
    .Q(\data_array.data1[4][38] ));
 sky130_fd_sc_hd__dfxtp_2 _13935_ (.CLK(clk),
    .D(_02564_),
    .Q(\data_array.data1[4][39] ));
 sky130_fd_sc_hd__dfxtp_2 _13936_ (.CLK(clk),
    .D(_02565_),
    .Q(\data_array.data1[4][40] ));
 sky130_fd_sc_hd__dfxtp_2 _13937_ (.CLK(clk),
    .D(_02566_),
    .Q(\data_array.data1[4][41] ));
 sky130_fd_sc_hd__dfxtp_2 _13938_ (.CLK(clk),
    .D(_02567_),
    .Q(\data_array.data1[4][42] ));
 sky130_fd_sc_hd__dfxtp_2 _13939_ (.CLK(clk),
    .D(_02568_),
    .Q(\data_array.data1[4][43] ));
 sky130_fd_sc_hd__dfxtp_2 _13940_ (.CLK(clk),
    .D(_02569_),
    .Q(\data_array.data1[4][44] ));
 sky130_fd_sc_hd__dfxtp_2 _13941_ (.CLK(clk),
    .D(_02570_),
    .Q(\data_array.data1[4][45] ));
 sky130_fd_sc_hd__dfxtp_2 _13942_ (.CLK(clk),
    .D(_02571_),
    .Q(\data_array.data1[4][46] ));
 sky130_fd_sc_hd__dfxtp_2 _13943_ (.CLK(clk),
    .D(_02572_),
    .Q(\data_array.data1[4][47] ));
 sky130_fd_sc_hd__dfxtp_2 _13944_ (.CLK(clk),
    .D(_02573_),
    .Q(\data_array.data1[4][48] ));
 sky130_fd_sc_hd__dfxtp_2 _13945_ (.CLK(clk),
    .D(_02574_),
    .Q(\data_array.data1[4][49] ));
 sky130_fd_sc_hd__dfxtp_2 _13946_ (.CLK(clk),
    .D(_02575_),
    .Q(\data_array.data1[4][50] ));
 sky130_fd_sc_hd__dfxtp_2 _13947_ (.CLK(clk),
    .D(_02576_),
    .Q(\data_array.data1[4][51] ));
 sky130_fd_sc_hd__dfxtp_2 _13948_ (.CLK(clk),
    .D(_02577_),
    .Q(\data_array.data1[4][52] ));
 sky130_fd_sc_hd__dfxtp_2 _13949_ (.CLK(clk),
    .D(_02578_),
    .Q(\data_array.data1[4][53] ));
 sky130_fd_sc_hd__dfxtp_2 _13950_ (.CLK(clk),
    .D(_02579_),
    .Q(\data_array.data1[4][54] ));
 sky130_fd_sc_hd__dfxtp_2 _13951_ (.CLK(clk),
    .D(_02580_),
    .Q(\data_array.data1[4][55] ));
 sky130_fd_sc_hd__dfxtp_2 _13952_ (.CLK(clk),
    .D(_02581_),
    .Q(\data_array.data1[4][56] ));
 sky130_fd_sc_hd__dfxtp_2 _13953_ (.CLK(clk),
    .D(_02582_),
    .Q(\data_array.data1[4][57] ));
 sky130_fd_sc_hd__dfxtp_2 _13954_ (.CLK(clk),
    .D(_02583_),
    .Q(\data_array.data1[4][58] ));
 sky130_fd_sc_hd__dfxtp_2 _13955_ (.CLK(clk),
    .D(_02584_),
    .Q(\data_array.data1[4][59] ));
 sky130_fd_sc_hd__dfxtp_2 _13956_ (.CLK(clk),
    .D(_02585_),
    .Q(\data_array.data1[4][60] ));
 sky130_fd_sc_hd__dfxtp_2 _13957_ (.CLK(clk),
    .D(_02586_),
    .Q(\data_array.data1[4][61] ));
 sky130_fd_sc_hd__dfxtp_2 _13958_ (.CLK(clk),
    .D(_02587_),
    .Q(\data_array.data1[4][62] ));
 sky130_fd_sc_hd__dfxtp_2 _13959_ (.CLK(clk),
    .D(_02588_),
    .Q(\data_array.data1[4][63] ));
 sky130_fd_sc_hd__dfxtp_2 _13960_ (.CLK(clk),
    .D(_02589_),
    .Q(\data_array.data1[5][0] ));
 sky130_fd_sc_hd__dfxtp_2 _13961_ (.CLK(clk),
    .D(_02590_),
    .Q(\data_array.data1[5][1] ));
 sky130_fd_sc_hd__dfxtp_2 _13962_ (.CLK(clk),
    .D(_02591_),
    .Q(\data_array.data1[5][2] ));
 sky130_fd_sc_hd__dfxtp_2 _13963_ (.CLK(clk),
    .D(_02592_),
    .Q(\data_array.data1[5][3] ));
 sky130_fd_sc_hd__dfxtp_2 _13964_ (.CLK(clk),
    .D(_02593_),
    .Q(\data_array.data1[5][4] ));
 sky130_fd_sc_hd__dfxtp_2 _13965_ (.CLK(clk),
    .D(_02594_),
    .Q(\data_array.data1[5][5] ));
 sky130_fd_sc_hd__dfxtp_2 _13966_ (.CLK(clk),
    .D(_02595_),
    .Q(\data_array.data1[5][6] ));
 sky130_fd_sc_hd__dfxtp_2 _13967_ (.CLK(clk),
    .D(_02596_),
    .Q(\data_array.data1[5][7] ));
 sky130_fd_sc_hd__dfxtp_2 _13968_ (.CLK(clk),
    .D(_02597_),
    .Q(\data_array.data1[5][8] ));
 sky130_fd_sc_hd__dfxtp_2 _13969_ (.CLK(clk),
    .D(_02598_),
    .Q(\data_array.data1[5][9] ));
 sky130_fd_sc_hd__dfxtp_2 _13970_ (.CLK(clk),
    .D(_02599_),
    .Q(\data_array.data1[5][10] ));
 sky130_fd_sc_hd__dfxtp_2 _13971_ (.CLK(clk),
    .D(_02600_),
    .Q(\data_array.data1[5][11] ));
 sky130_fd_sc_hd__dfxtp_2 _13972_ (.CLK(clk),
    .D(_02601_),
    .Q(\data_array.data1[5][12] ));
 sky130_fd_sc_hd__dfxtp_2 _13973_ (.CLK(clk),
    .D(_02602_),
    .Q(\data_array.data1[5][13] ));
 sky130_fd_sc_hd__dfxtp_2 _13974_ (.CLK(clk),
    .D(_02603_),
    .Q(\data_array.data1[5][14] ));
 sky130_fd_sc_hd__dfxtp_2 _13975_ (.CLK(clk),
    .D(_02604_),
    .Q(\data_array.data1[5][15] ));
 sky130_fd_sc_hd__dfxtp_2 _13976_ (.CLK(clk),
    .D(_02605_),
    .Q(\data_array.data1[5][16] ));
 sky130_fd_sc_hd__dfxtp_2 _13977_ (.CLK(clk),
    .D(_02606_),
    .Q(\data_array.data1[5][17] ));
 sky130_fd_sc_hd__dfxtp_2 _13978_ (.CLK(clk),
    .D(_02607_),
    .Q(\data_array.data1[5][18] ));
 sky130_fd_sc_hd__dfxtp_2 _13979_ (.CLK(clk),
    .D(_02608_),
    .Q(\data_array.data1[5][19] ));
 sky130_fd_sc_hd__dfxtp_2 _13980_ (.CLK(clk),
    .D(_02609_),
    .Q(\data_array.data1[5][20] ));
 sky130_fd_sc_hd__dfxtp_2 _13981_ (.CLK(clk),
    .D(_02610_),
    .Q(\data_array.data1[5][21] ));
 sky130_fd_sc_hd__dfxtp_2 _13982_ (.CLK(clk),
    .D(_02611_),
    .Q(\data_array.data1[5][22] ));
 sky130_fd_sc_hd__dfxtp_2 _13983_ (.CLK(clk),
    .D(_02612_),
    .Q(\data_array.data1[5][23] ));
 sky130_fd_sc_hd__dfxtp_2 _13984_ (.CLK(clk),
    .D(_02613_),
    .Q(\data_array.data1[5][24] ));
 sky130_fd_sc_hd__dfxtp_2 _13985_ (.CLK(clk),
    .D(_02614_),
    .Q(\data_array.data1[5][25] ));
 sky130_fd_sc_hd__dfxtp_2 _13986_ (.CLK(clk),
    .D(_02615_),
    .Q(\data_array.data1[5][26] ));
 sky130_fd_sc_hd__dfxtp_2 _13987_ (.CLK(clk),
    .D(_02616_),
    .Q(\data_array.data1[5][27] ));
 sky130_fd_sc_hd__dfxtp_2 _13988_ (.CLK(clk),
    .D(_02617_),
    .Q(\data_array.data1[5][28] ));
 sky130_fd_sc_hd__dfxtp_2 _13989_ (.CLK(clk),
    .D(_02618_),
    .Q(\data_array.data1[5][29] ));
 sky130_fd_sc_hd__dfxtp_2 _13990_ (.CLK(clk),
    .D(_02619_),
    .Q(\data_array.data1[5][30] ));
 sky130_fd_sc_hd__dfxtp_2 _13991_ (.CLK(clk),
    .D(_02620_),
    .Q(\data_array.data1[5][31] ));
 sky130_fd_sc_hd__dfxtp_2 _13992_ (.CLK(clk),
    .D(_02621_),
    .Q(\data_array.data1[5][32] ));
 sky130_fd_sc_hd__dfxtp_2 _13993_ (.CLK(clk),
    .D(_02622_),
    .Q(\data_array.data1[5][33] ));
 sky130_fd_sc_hd__dfxtp_2 _13994_ (.CLK(clk),
    .D(_02623_),
    .Q(\data_array.data1[5][34] ));
 sky130_fd_sc_hd__dfxtp_2 _13995_ (.CLK(clk),
    .D(_02624_),
    .Q(\data_array.data1[5][35] ));
 sky130_fd_sc_hd__dfxtp_2 _13996_ (.CLK(clk),
    .D(_02625_),
    .Q(\data_array.data1[5][36] ));
 sky130_fd_sc_hd__dfxtp_2 _13997_ (.CLK(clk),
    .D(_02626_),
    .Q(\data_array.data1[5][37] ));
 sky130_fd_sc_hd__dfxtp_2 _13998_ (.CLK(clk),
    .D(_02627_),
    .Q(\data_array.data1[5][38] ));
 sky130_fd_sc_hd__dfxtp_2 _13999_ (.CLK(clk),
    .D(_02628_),
    .Q(\data_array.data1[5][39] ));
 sky130_fd_sc_hd__dfxtp_2 _14000_ (.CLK(clk),
    .D(_02629_),
    .Q(\data_array.data1[5][40] ));
 sky130_fd_sc_hd__dfxtp_2 _14001_ (.CLK(clk),
    .D(_02630_),
    .Q(\data_array.data1[5][41] ));
 sky130_fd_sc_hd__dfxtp_2 _14002_ (.CLK(clk),
    .D(_02631_),
    .Q(\data_array.data1[5][42] ));
 sky130_fd_sc_hd__dfxtp_2 _14003_ (.CLK(clk),
    .D(_02632_),
    .Q(\data_array.data1[5][43] ));
 sky130_fd_sc_hd__dfxtp_2 _14004_ (.CLK(clk),
    .D(_02633_),
    .Q(\data_array.data1[5][44] ));
 sky130_fd_sc_hd__dfxtp_2 _14005_ (.CLK(clk),
    .D(_02634_),
    .Q(\data_array.data1[5][45] ));
 sky130_fd_sc_hd__dfxtp_2 _14006_ (.CLK(clk),
    .D(_02635_),
    .Q(\data_array.data1[5][46] ));
 sky130_fd_sc_hd__dfxtp_2 _14007_ (.CLK(clk),
    .D(_02636_),
    .Q(\data_array.data1[5][47] ));
 sky130_fd_sc_hd__dfxtp_2 _14008_ (.CLK(clk),
    .D(_02637_),
    .Q(\data_array.data1[5][48] ));
 sky130_fd_sc_hd__dfxtp_2 _14009_ (.CLK(clk),
    .D(_02638_),
    .Q(\data_array.data1[5][49] ));
 sky130_fd_sc_hd__dfxtp_2 _14010_ (.CLK(clk),
    .D(_02639_),
    .Q(\data_array.data1[5][50] ));
 sky130_fd_sc_hd__dfxtp_2 _14011_ (.CLK(clk),
    .D(_02640_),
    .Q(\data_array.data1[5][51] ));
 sky130_fd_sc_hd__dfxtp_2 _14012_ (.CLK(clk),
    .D(_02641_),
    .Q(\data_array.data1[5][52] ));
 sky130_fd_sc_hd__dfxtp_2 _14013_ (.CLK(clk),
    .D(_02642_),
    .Q(\data_array.data1[5][53] ));
 sky130_fd_sc_hd__dfxtp_2 _14014_ (.CLK(clk),
    .D(_02643_),
    .Q(\data_array.data1[5][54] ));
 sky130_fd_sc_hd__dfxtp_2 _14015_ (.CLK(clk),
    .D(_02644_),
    .Q(\data_array.data1[5][55] ));
 sky130_fd_sc_hd__dfxtp_2 _14016_ (.CLK(clk),
    .D(_02645_),
    .Q(\data_array.data1[5][56] ));
 sky130_fd_sc_hd__dfxtp_2 _14017_ (.CLK(clk),
    .D(_02646_),
    .Q(\data_array.data1[5][57] ));
 sky130_fd_sc_hd__dfxtp_2 _14018_ (.CLK(clk),
    .D(_02647_),
    .Q(\data_array.data1[5][58] ));
 sky130_fd_sc_hd__dfxtp_2 _14019_ (.CLK(clk),
    .D(_02648_),
    .Q(\data_array.data1[5][59] ));
 sky130_fd_sc_hd__dfxtp_2 _14020_ (.CLK(clk),
    .D(_02649_),
    .Q(\data_array.data1[5][60] ));
 sky130_fd_sc_hd__dfxtp_2 _14021_ (.CLK(clk),
    .D(_02650_),
    .Q(\data_array.data1[5][61] ));
 sky130_fd_sc_hd__dfxtp_2 _14022_ (.CLK(clk),
    .D(_02651_),
    .Q(\data_array.data1[5][62] ));
 sky130_fd_sc_hd__dfxtp_2 _14023_ (.CLK(clk),
    .D(_02652_),
    .Q(\data_array.data1[5][63] ));
 sky130_fd_sc_hd__dfxtp_2 _14024_ (.CLK(clk),
    .D(_02653_),
    .Q(\data_array.data1[6][0] ));
 sky130_fd_sc_hd__dfxtp_2 _14025_ (.CLK(clk),
    .D(_02654_),
    .Q(\data_array.data1[6][1] ));
 sky130_fd_sc_hd__dfxtp_2 _14026_ (.CLK(clk),
    .D(_02655_),
    .Q(\data_array.data1[6][2] ));
 sky130_fd_sc_hd__dfxtp_2 _14027_ (.CLK(clk),
    .D(_02656_),
    .Q(\data_array.data1[6][3] ));
 sky130_fd_sc_hd__dfxtp_2 _14028_ (.CLK(clk),
    .D(_02657_),
    .Q(\data_array.data1[6][4] ));
 sky130_fd_sc_hd__dfxtp_2 _14029_ (.CLK(clk),
    .D(_02658_),
    .Q(\data_array.data1[6][5] ));
 sky130_fd_sc_hd__dfxtp_2 _14030_ (.CLK(clk),
    .D(_02659_),
    .Q(\data_array.data1[6][6] ));
 sky130_fd_sc_hd__dfxtp_2 _14031_ (.CLK(clk),
    .D(_02660_),
    .Q(\data_array.data1[6][7] ));
 sky130_fd_sc_hd__dfxtp_2 _14032_ (.CLK(clk),
    .D(_02661_),
    .Q(\data_array.data1[6][8] ));
 sky130_fd_sc_hd__dfxtp_2 _14033_ (.CLK(clk),
    .D(_02662_),
    .Q(\data_array.data1[6][9] ));
 sky130_fd_sc_hd__dfxtp_2 _14034_ (.CLK(clk),
    .D(_02663_),
    .Q(\data_array.data1[6][10] ));
 sky130_fd_sc_hd__dfxtp_2 _14035_ (.CLK(clk),
    .D(_02664_),
    .Q(\data_array.data1[6][11] ));
 sky130_fd_sc_hd__dfxtp_2 _14036_ (.CLK(clk),
    .D(_02665_),
    .Q(\data_array.data1[6][12] ));
 sky130_fd_sc_hd__dfxtp_2 _14037_ (.CLK(clk),
    .D(_02666_),
    .Q(\data_array.data1[6][13] ));
 sky130_fd_sc_hd__dfxtp_2 _14038_ (.CLK(clk),
    .D(_02667_),
    .Q(\data_array.data1[6][14] ));
 sky130_fd_sc_hd__dfxtp_2 _14039_ (.CLK(clk),
    .D(_02668_),
    .Q(\data_array.data1[6][15] ));
 sky130_fd_sc_hd__dfxtp_2 _14040_ (.CLK(clk),
    .D(_02669_),
    .Q(\data_array.data1[6][16] ));
 sky130_fd_sc_hd__dfxtp_2 _14041_ (.CLK(clk),
    .D(_02670_),
    .Q(\data_array.data1[6][17] ));
 sky130_fd_sc_hd__dfxtp_2 _14042_ (.CLK(clk),
    .D(_02671_),
    .Q(\data_array.data1[6][18] ));
 sky130_fd_sc_hd__dfxtp_2 _14043_ (.CLK(clk),
    .D(_02672_),
    .Q(\data_array.data1[6][19] ));
 sky130_fd_sc_hd__dfxtp_2 _14044_ (.CLK(clk),
    .D(_02673_),
    .Q(\data_array.data1[6][20] ));
 sky130_fd_sc_hd__dfxtp_2 _14045_ (.CLK(clk),
    .D(_02674_),
    .Q(\data_array.data1[6][21] ));
 sky130_fd_sc_hd__dfxtp_2 _14046_ (.CLK(clk),
    .D(_02675_),
    .Q(\data_array.data1[6][22] ));
 sky130_fd_sc_hd__dfxtp_2 _14047_ (.CLK(clk),
    .D(_02676_),
    .Q(\data_array.data1[6][23] ));
 sky130_fd_sc_hd__dfxtp_2 _14048_ (.CLK(clk),
    .D(_02677_),
    .Q(\data_array.data1[6][24] ));
 sky130_fd_sc_hd__dfxtp_2 _14049_ (.CLK(clk),
    .D(_02678_),
    .Q(\data_array.data1[6][25] ));
 sky130_fd_sc_hd__dfxtp_2 _14050_ (.CLK(clk),
    .D(_02679_),
    .Q(\data_array.data1[6][26] ));
 sky130_fd_sc_hd__dfxtp_2 _14051_ (.CLK(clk),
    .D(_02680_),
    .Q(\data_array.data1[6][27] ));
 sky130_fd_sc_hd__dfxtp_2 _14052_ (.CLK(clk),
    .D(_02681_),
    .Q(\data_array.data1[6][28] ));
 sky130_fd_sc_hd__dfxtp_2 _14053_ (.CLK(clk),
    .D(_02682_),
    .Q(\data_array.data1[6][29] ));
 sky130_fd_sc_hd__dfxtp_2 _14054_ (.CLK(clk),
    .D(_02683_),
    .Q(\data_array.data1[6][30] ));
 sky130_fd_sc_hd__dfxtp_2 _14055_ (.CLK(clk),
    .D(_02684_),
    .Q(\data_array.data1[6][31] ));
 sky130_fd_sc_hd__dfxtp_2 _14056_ (.CLK(clk),
    .D(_02685_),
    .Q(\data_array.data1[6][32] ));
 sky130_fd_sc_hd__dfxtp_2 _14057_ (.CLK(clk),
    .D(_02686_),
    .Q(\data_array.data1[6][33] ));
 sky130_fd_sc_hd__dfxtp_2 _14058_ (.CLK(clk),
    .D(_02687_),
    .Q(\data_array.data1[6][34] ));
 sky130_fd_sc_hd__dfxtp_2 _14059_ (.CLK(clk),
    .D(_02688_),
    .Q(\data_array.data1[6][35] ));
 sky130_fd_sc_hd__dfxtp_2 _14060_ (.CLK(clk),
    .D(_02689_),
    .Q(\data_array.data1[6][36] ));
 sky130_fd_sc_hd__dfxtp_2 _14061_ (.CLK(clk),
    .D(_02690_),
    .Q(\data_array.data1[6][37] ));
 sky130_fd_sc_hd__dfxtp_2 _14062_ (.CLK(clk),
    .D(_02691_),
    .Q(\data_array.data1[6][38] ));
 sky130_fd_sc_hd__dfxtp_2 _14063_ (.CLK(clk),
    .D(_02692_),
    .Q(\data_array.data1[6][39] ));
 sky130_fd_sc_hd__dfxtp_2 _14064_ (.CLK(clk),
    .D(_02693_),
    .Q(\data_array.data1[6][40] ));
 sky130_fd_sc_hd__dfxtp_2 _14065_ (.CLK(clk),
    .D(_02694_),
    .Q(\data_array.data1[6][41] ));
 sky130_fd_sc_hd__dfxtp_2 _14066_ (.CLK(clk),
    .D(_02695_),
    .Q(\data_array.data1[6][42] ));
 sky130_fd_sc_hd__dfxtp_2 _14067_ (.CLK(clk),
    .D(_02696_),
    .Q(\data_array.data1[6][43] ));
 sky130_fd_sc_hd__dfxtp_2 _14068_ (.CLK(clk),
    .D(_02697_),
    .Q(\data_array.data1[6][44] ));
 sky130_fd_sc_hd__dfxtp_2 _14069_ (.CLK(clk),
    .D(_02698_),
    .Q(\data_array.data1[6][45] ));
 sky130_fd_sc_hd__dfxtp_2 _14070_ (.CLK(clk),
    .D(_02699_),
    .Q(\data_array.data1[6][46] ));
 sky130_fd_sc_hd__dfxtp_2 _14071_ (.CLK(clk),
    .D(_02700_),
    .Q(\data_array.data1[6][47] ));
 sky130_fd_sc_hd__dfxtp_2 _14072_ (.CLK(clk),
    .D(_02701_),
    .Q(\data_array.data1[6][48] ));
 sky130_fd_sc_hd__dfxtp_2 _14073_ (.CLK(clk),
    .D(_02702_),
    .Q(\data_array.data1[6][49] ));
 sky130_fd_sc_hd__dfxtp_2 _14074_ (.CLK(clk),
    .D(_02703_),
    .Q(\data_array.data1[6][50] ));
 sky130_fd_sc_hd__dfxtp_2 _14075_ (.CLK(clk),
    .D(_02704_),
    .Q(\data_array.data1[6][51] ));
 sky130_fd_sc_hd__dfxtp_2 _14076_ (.CLK(clk),
    .D(_02705_),
    .Q(\data_array.data1[6][52] ));
 sky130_fd_sc_hd__dfxtp_2 _14077_ (.CLK(clk),
    .D(_02706_),
    .Q(\data_array.data1[6][53] ));
 sky130_fd_sc_hd__dfxtp_2 _14078_ (.CLK(clk),
    .D(_02707_),
    .Q(\data_array.data1[6][54] ));
 sky130_fd_sc_hd__dfxtp_2 _14079_ (.CLK(clk),
    .D(_02708_),
    .Q(\data_array.data1[6][55] ));
 sky130_fd_sc_hd__dfxtp_2 _14080_ (.CLK(clk),
    .D(_02709_),
    .Q(\data_array.data1[6][56] ));
 sky130_fd_sc_hd__dfxtp_2 _14081_ (.CLK(clk),
    .D(_02710_),
    .Q(\data_array.data1[6][57] ));
 sky130_fd_sc_hd__dfxtp_2 _14082_ (.CLK(clk),
    .D(_02711_),
    .Q(\data_array.data1[6][58] ));
 sky130_fd_sc_hd__dfxtp_2 _14083_ (.CLK(clk),
    .D(_02712_),
    .Q(\data_array.data1[6][59] ));
 sky130_fd_sc_hd__dfxtp_2 _14084_ (.CLK(clk),
    .D(_02713_),
    .Q(\data_array.data1[6][60] ));
 sky130_fd_sc_hd__dfxtp_2 _14085_ (.CLK(clk),
    .D(_02714_),
    .Q(\data_array.data1[6][61] ));
 sky130_fd_sc_hd__dfxtp_2 _14086_ (.CLK(clk),
    .D(_02715_),
    .Q(\data_array.data1[6][62] ));
 sky130_fd_sc_hd__dfxtp_2 _14087_ (.CLK(clk),
    .D(_02716_),
    .Q(\data_array.data1[6][63] ));
 sky130_fd_sc_hd__dfxtp_2 _14088_ (.CLK(clk),
    .D(_02717_),
    .Q(\data_array.data0[1][0] ));
 sky130_fd_sc_hd__dfxtp_2 _14089_ (.CLK(clk),
    .D(_02718_),
    .Q(\data_array.data0[1][1] ));
 sky130_fd_sc_hd__dfxtp_2 _14090_ (.CLK(clk),
    .D(_02719_),
    .Q(\data_array.data0[1][2] ));
 sky130_fd_sc_hd__dfxtp_2 _14091_ (.CLK(clk),
    .D(_02720_),
    .Q(\data_array.data0[1][3] ));
 sky130_fd_sc_hd__dfxtp_2 _14092_ (.CLK(clk),
    .D(_02721_),
    .Q(\data_array.data0[1][4] ));
 sky130_fd_sc_hd__dfxtp_2 _14093_ (.CLK(clk),
    .D(_02722_),
    .Q(\data_array.data0[1][5] ));
 sky130_fd_sc_hd__dfxtp_2 _14094_ (.CLK(clk),
    .D(_02723_),
    .Q(\data_array.data0[1][6] ));
 sky130_fd_sc_hd__dfxtp_2 _14095_ (.CLK(clk),
    .D(_02724_),
    .Q(\data_array.data0[1][7] ));
 sky130_fd_sc_hd__dfxtp_2 _14096_ (.CLK(clk),
    .D(_02725_),
    .Q(\data_array.data0[1][8] ));
 sky130_fd_sc_hd__dfxtp_2 _14097_ (.CLK(clk),
    .D(_02726_),
    .Q(\data_array.data0[1][9] ));
 sky130_fd_sc_hd__dfxtp_2 _14098_ (.CLK(clk),
    .D(_02727_),
    .Q(\data_array.data0[1][10] ));
 sky130_fd_sc_hd__dfxtp_2 _14099_ (.CLK(clk),
    .D(_02728_),
    .Q(\data_array.data0[1][11] ));
 sky130_fd_sc_hd__dfxtp_2 _14100_ (.CLK(clk),
    .D(_02729_),
    .Q(\data_array.data0[1][12] ));
 sky130_fd_sc_hd__dfxtp_2 _14101_ (.CLK(clk),
    .D(_02730_),
    .Q(\data_array.data0[1][13] ));
 sky130_fd_sc_hd__dfxtp_2 _14102_ (.CLK(clk),
    .D(_02731_),
    .Q(\data_array.data0[1][14] ));
 sky130_fd_sc_hd__dfxtp_2 _14103_ (.CLK(clk),
    .D(_02732_),
    .Q(\data_array.data0[1][15] ));
 sky130_fd_sc_hd__dfxtp_2 _14104_ (.CLK(clk),
    .D(_02733_),
    .Q(\data_array.data0[1][16] ));
 sky130_fd_sc_hd__dfxtp_2 _14105_ (.CLK(clk),
    .D(_02734_),
    .Q(\data_array.data0[1][17] ));
 sky130_fd_sc_hd__dfxtp_2 _14106_ (.CLK(clk),
    .D(_02735_),
    .Q(\data_array.data0[1][18] ));
 sky130_fd_sc_hd__dfxtp_2 _14107_ (.CLK(clk),
    .D(_02736_),
    .Q(\data_array.data0[1][19] ));
 sky130_fd_sc_hd__dfxtp_2 _14108_ (.CLK(clk),
    .D(_02737_),
    .Q(\data_array.data0[1][20] ));
 sky130_fd_sc_hd__dfxtp_2 _14109_ (.CLK(clk),
    .D(_02738_),
    .Q(\data_array.data0[1][21] ));
 sky130_fd_sc_hd__dfxtp_2 _14110_ (.CLK(clk),
    .D(_02739_),
    .Q(\data_array.data0[1][22] ));
 sky130_fd_sc_hd__dfxtp_2 _14111_ (.CLK(clk),
    .D(_02740_),
    .Q(\data_array.data0[1][23] ));
 sky130_fd_sc_hd__dfxtp_2 _14112_ (.CLK(clk),
    .D(_02741_),
    .Q(\data_array.data0[1][24] ));
 sky130_fd_sc_hd__dfxtp_2 _14113_ (.CLK(clk),
    .D(_02742_),
    .Q(\data_array.data0[1][25] ));
 sky130_fd_sc_hd__dfxtp_2 _14114_ (.CLK(clk),
    .D(_02743_),
    .Q(\data_array.data0[1][26] ));
 sky130_fd_sc_hd__dfxtp_2 _14115_ (.CLK(clk),
    .D(_02744_),
    .Q(\data_array.data0[1][27] ));
 sky130_fd_sc_hd__dfxtp_2 _14116_ (.CLK(clk),
    .D(_02745_),
    .Q(\data_array.data0[1][28] ));
 sky130_fd_sc_hd__dfxtp_2 _14117_ (.CLK(clk),
    .D(_02746_),
    .Q(\data_array.data0[1][29] ));
 sky130_fd_sc_hd__dfxtp_2 _14118_ (.CLK(clk),
    .D(_02747_),
    .Q(\data_array.data0[1][30] ));
 sky130_fd_sc_hd__dfxtp_2 _14119_ (.CLK(clk),
    .D(_02748_),
    .Q(\data_array.data0[1][31] ));
 sky130_fd_sc_hd__dfxtp_2 _14120_ (.CLK(clk),
    .D(_02749_),
    .Q(\data_array.data0[1][32] ));
 sky130_fd_sc_hd__dfxtp_2 _14121_ (.CLK(clk),
    .D(_02750_),
    .Q(\data_array.data0[1][33] ));
 sky130_fd_sc_hd__dfxtp_2 _14122_ (.CLK(clk),
    .D(_02751_),
    .Q(\data_array.data0[1][34] ));
 sky130_fd_sc_hd__dfxtp_2 _14123_ (.CLK(clk),
    .D(_02752_),
    .Q(\data_array.data0[1][35] ));
 sky130_fd_sc_hd__dfxtp_2 _14124_ (.CLK(clk),
    .D(_02753_),
    .Q(\data_array.data0[1][36] ));
 sky130_fd_sc_hd__dfxtp_2 _14125_ (.CLK(clk),
    .D(_02754_),
    .Q(\data_array.data0[1][37] ));
 sky130_fd_sc_hd__dfxtp_2 _14126_ (.CLK(clk),
    .D(_02755_),
    .Q(\data_array.data0[1][38] ));
 sky130_fd_sc_hd__dfxtp_2 _14127_ (.CLK(clk),
    .D(_02756_),
    .Q(\data_array.data0[1][39] ));
 sky130_fd_sc_hd__dfxtp_2 _14128_ (.CLK(clk),
    .D(_02757_),
    .Q(\data_array.data0[1][40] ));
 sky130_fd_sc_hd__dfxtp_2 _14129_ (.CLK(clk),
    .D(_02758_),
    .Q(\data_array.data0[1][41] ));
 sky130_fd_sc_hd__dfxtp_2 _14130_ (.CLK(clk),
    .D(_02759_),
    .Q(\data_array.data0[1][42] ));
 sky130_fd_sc_hd__dfxtp_2 _14131_ (.CLK(clk),
    .D(_02760_),
    .Q(\data_array.data0[1][43] ));
 sky130_fd_sc_hd__dfxtp_2 _14132_ (.CLK(clk),
    .D(_02761_),
    .Q(\data_array.data0[1][44] ));
 sky130_fd_sc_hd__dfxtp_2 _14133_ (.CLK(clk),
    .D(_02762_),
    .Q(\data_array.data0[1][45] ));
 sky130_fd_sc_hd__dfxtp_2 _14134_ (.CLK(clk),
    .D(_02763_),
    .Q(\data_array.data0[1][46] ));
 sky130_fd_sc_hd__dfxtp_2 _14135_ (.CLK(clk),
    .D(_02764_),
    .Q(\data_array.data0[1][47] ));
 sky130_fd_sc_hd__dfxtp_2 _14136_ (.CLK(clk),
    .D(_02765_),
    .Q(\data_array.data0[1][48] ));
 sky130_fd_sc_hd__dfxtp_2 _14137_ (.CLK(clk),
    .D(_02766_),
    .Q(\data_array.data0[1][49] ));
 sky130_fd_sc_hd__dfxtp_2 _14138_ (.CLK(clk),
    .D(_02767_),
    .Q(\data_array.data0[1][50] ));
 sky130_fd_sc_hd__dfxtp_2 _14139_ (.CLK(clk),
    .D(_02768_),
    .Q(\data_array.data0[1][51] ));
 sky130_fd_sc_hd__dfxtp_2 _14140_ (.CLK(clk),
    .D(_02769_),
    .Q(\data_array.data0[1][52] ));
 sky130_fd_sc_hd__dfxtp_2 _14141_ (.CLK(clk),
    .D(_02770_),
    .Q(\data_array.data0[1][53] ));
 sky130_fd_sc_hd__dfxtp_2 _14142_ (.CLK(clk),
    .D(_02771_),
    .Q(\data_array.data0[1][54] ));
 sky130_fd_sc_hd__dfxtp_2 _14143_ (.CLK(clk),
    .D(_02772_),
    .Q(\data_array.data0[1][55] ));
 sky130_fd_sc_hd__dfxtp_2 _14144_ (.CLK(clk),
    .D(_02773_),
    .Q(\data_array.data0[1][56] ));
 sky130_fd_sc_hd__dfxtp_2 _14145_ (.CLK(clk),
    .D(_02774_),
    .Q(\data_array.data0[1][57] ));
 sky130_fd_sc_hd__dfxtp_2 _14146_ (.CLK(clk),
    .D(_02775_),
    .Q(\data_array.data0[1][58] ));
 sky130_fd_sc_hd__dfxtp_2 _14147_ (.CLK(clk),
    .D(_02776_),
    .Q(\data_array.data0[1][59] ));
 sky130_fd_sc_hd__dfxtp_2 _14148_ (.CLK(clk),
    .D(_02777_),
    .Q(\data_array.data0[1][60] ));
 sky130_fd_sc_hd__dfxtp_2 _14149_ (.CLK(clk),
    .D(_02778_),
    .Q(\data_array.data0[1][61] ));
 sky130_fd_sc_hd__dfxtp_2 _14150_ (.CLK(clk),
    .D(_02779_),
    .Q(\data_array.data0[1][62] ));
 sky130_fd_sc_hd__dfxtp_2 _14151_ (.CLK(clk),
    .D(_02780_),
    .Q(\data_array.data0[1][63] ));
 sky130_fd_sc_hd__dfxtp_2 _14152_ (.CLK(clk),
    .D(_02781_),
    .Q(\data_array.data0[2][0] ));
 sky130_fd_sc_hd__dfxtp_2 _14153_ (.CLK(clk),
    .D(_02782_),
    .Q(\data_array.data0[2][1] ));
 sky130_fd_sc_hd__dfxtp_2 _14154_ (.CLK(clk),
    .D(_02783_),
    .Q(\data_array.data0[2][2] ));
 sky130_fd_sc_hd__dfxtp_2 _14155_ (.CLK(clk),
    .D(_02784_),
    .Q(\data_array.data0[2][3] ));
 sky130_fd_sc_hd__dfxtp_2 _14156_ (.CLK(clk),
    .D(_02785_),
    .Q(\data_array.data0[2][4] ));
 sky130_fd_sc_hd__dfxtp_2 _14157_ (.CLK(clk),
    .D(_02786_),
    .Q(\data_array.data0[2][5] ));
 sky130_fd_sc_hd__dfxtp_2 _14158_ (.CLK(clk),
    .D(_02787_),
    .Q(\data_array.data0[2][6] ));
 sky130_fd_sc_hd__dfxtp_2 _14159_ (.CLK(clk),
    .D(_02788_),
    .Q(\data_array.data0[2][7] ));
 sky130_fd_sc_hd__dfxtp_2 _14160_ (.CLK(clk),
    .D(_02789_),
    .Q(\data_array.data0[2][8] ));
 sky130_fd_sc_hd__dfxtp_2 _14161_ (.CLK(clk),
    .D(_02790_),
    .Q(\data_array.data0[2][9] ));
 sky130_fd_sc_hd__dfxtp_2 _14162_ (.CLK(clk),
    .D(_02791_),
    .Q(\data_array.data0[2][10] ));
 sky130_fd_sc_hd__dfxtp_2 _14163_ (.CLK(clk),
    .D(_02792_),
    .Q(\data_array.data0[2][11] ));
 sky130_fd_sc_hd__dfxtp_2 _14164_ (.CLK(clk),
    .D(_02793_),
    .Q(\data_array.data0[2][12] ));
 sky130_fd_sc_hd__dfxtp_2 _14165_ (.CLK(clk),
    .D(_02794_),
    .Q(\data_array.data0[2][13] ));
 sky130_fd_sc_hd__dfxtp_2 _14166_ (.CLK(clk),
    .D(_02795_),
    .Q(\data_array.data0[2][14] ));
 sky130_fd_sc_hd__dfxtp_2 _14167_ (.CLK(clk),
    .D(_02796_),
    .Q(\data_array.data0[2][15] ));
 sky130_fd_sc_hd__dfxtp_2 _14168_ (.CLK(clk),
    .D(_02797_),
    .Q(\data_array.data0[2][16] ));
 sky130_fd_sc_hd__dfxtp_2 _14169_ (.CLK(clk),
    .D(_02798_),
    .Q(\data_array.data0[2][17] ));
 sky130_fd_sc_hd__dfxtp_2 _14170_ (.CLK(clk),
    .D(_02799_),
    .Q(\data_array.data0[2][18] ));
 sky130_fd_sc_hd__dfxtp_2 _14171_ (.CLK(clk),
    .D(_02800_),
    .Q(\data_array.data0[2][19] ));
 sky130_fd_sc_hd__dfxtp_2 _14172_ (.CLK(clk),
    .D(_02801_),
    .Q(\data_array.data0[2][20] ));
 sky130_fd_sc_hd__dfxtp_2 _14173_ (.CLK(clk),
    .D(_02802_),
    .Q(\data_array.data0[2][21] ));
 sky130_fd_sc_hd__dfxtp_2 _14174_ (.CLK(clk),
    .D(_02803_),
    .Q(\data_array.data0[2][22] ));
 sky130_fd_sc_hd__dfxtp_2 _14175_ (.CLK(clk),
    .D(_02804_),
    .Q(\data_array.data0[2][23] ));
 sky130_fd_sc_hd__dfxtp_2 _14176_ (.CLK(clk),
    .D(_02805_),
    .Q(\data_array.data0[2][24] ));
 sky130_fd_sc_hd__dfxtp_2 _14177_ (.CLK(clk),
    .D(_02806_),
    .Q(\data_array.data0[2][25] ));
 sky130_fd_sc_hd__dfxtp_2 _14178_ (.CLK(clk),
    .D(_02807_),
    .Q(\data_array.data0[2][26] ));
 sky130_fd_sc_hd__dfxtp_2 _14179_ (.CLK(clk),
    .D(_02808_),
    .Q(\data_array.data0[2][27] ));
 sky130_fd_sc_hd__dfxtp_2 _14180_ (.CLK(clk),
    .D(_02809_),
    .Q(\data_array.data0[2][28] ));
 sky130_fd_sc_hd__dfxtp_2 _14181_ (.CLK(clk),
    .D(_02810_),
    .Q(\data_array.data0[2][29] ));
 sky130_fd_sc_hd__dfxtp_2 _14182_ (.CLK(clk),
    .D(_02811_),
    .Q(\data_array.data0[2][30] ));
 sky130_fd_sc_hd__dfxtp_2 _14183_ (.CLK(clk),
    .D(_02812_),
    .Q(\data_array.data0[2][31] ));
 sky130_fd_sc_hd__dfxtp_2 _14184_ (.CLK(clk),
    .D(_02813_),
    .Q(\data_array.data0[2][32] ));
 sky130_fd_sc_hd__dfxtp_2 _14185_ (.CLK(clk),
    .D(_02814_),
    .Q(\data_array.data0[2][33] ));
 sky130_fd_sc_hd__dfxtp_2 _14186_ (.CLK(clk),
    .D(_02815_),
    .Q(\data_array.data0[2][34] ));
 sky130_fd_sc_hd__dfxtp_2 _14187_ (.CLK(clk),
    .D(_02816_),
    .Q(\data_array.data0[2][35] ));
 sky130_fd_sc_hd__dfxtp_2 _14188_ (.CLK(clk),
    .D(_02817_),
    .Q(\data_array.data0[2][36] ));
 sky130_fd_sc_hd__dfxtp_2 _14189_ (.CLK(clk),
    .D(_02818_),
    .Q(\data_array.data0[2][37] ));
 sky130_fd_sc_hd__dfxtp_2 _14190_ (.CLK(clk),
    .D(_02819_),
    .Q(\data_array.data0[2][38] ));
 sky130_fd_sc_hd__dfxtp_2 _14191_ (.CLK(clk),
    .D(_02820_),
    .Q(\data_array.data0[2][39] ));
 sky130_fd_sc_hd__dfxtp_2 _14192_ (.CLK(clk),
    .D(_02821_),
    .Q(\data_array.data0[2][40] ));
 sky130_fd_sc_hd__dfxtp_2 _14193_ (.CLK(clk),
    .D(_02822_),
    .Q(\data_array.data0[2][41] ));
 sky130_fd_sc_hd__dfxtp_2 _14194_ (.CLK(clk),
    .D(_02823_),
    .Q(\data_array.data0[2][42] ));
 sky130_fd_sc_hd__dfxtp_2 _14195_ (.CLK(clk),
    .D(_02824_),
    .Q(\data_array.data0[2][43] ));
 sky130_fd_sc_hd__dfxtp_2 _14196_ (.CLK(clk),
    .D(_02825_),
    .Q(\data_array.data0[2][44] ));
 sky130_fd_sc_hd__dfxtp_2 _14197_ (.CLK(clk),
    .D(_02826_),
    .Q(\data_array.data0[2][45] ));
 sky130_fd_sc_hd__dfxtp_2 _14198_ (.CLK(clk),
    .D(_02827_),
    .Q(\data_array.data0[2][46] ));
 sky130_fd_sc_hd__dfxtp_2 _14199_ (.CLK(clk),
    .D(_02828_),
    .Q(\data_array.data0[2][47] ));
 sky130_fd_sc_hd__dfxtp_2 _14200_ (.CLK(clk),
    .D(_02829_),
    .Q(\data_array.data0[2][48] ));
 sky130_fd_sc_hd__dfxtp_2 _14201_ (.CLK(clk),
    .D(_02830_),
    .Q(\data_array.data0[2][49] ));
 sky130_fd_sc_hd__dfxtp_2 _14202_ (.CLK(clk),
    .D(_02831_),
    .Q(\data_array.data0[2][50] ));
 sky130_fd_sc_hd__dfxtp_2 _14203_ (.CLK(clk),
    .D(_02832_),
    .Q(\data_array.data0[2][51] ));
 sky130_fd_sc_hd__dfxtp_2 _14204_ (.CLK(clk),
    .D(_02833_),
    .Q(\data_array.data0[2][52] ));
 sky130_fd_sc_hd__dfxtp_2 _14205_ (.CLK(clk),
    .D(_02834_),
    .Q(\data_array.data0[2][53] ));
 sky130_fd_sc_hd__dfxtp_2 _14206_ (.CLK(clk),
    .D(_02835_),
    .Q(\data_array.data0[2][54] ));
 sky130_fd_sc_hd__dfxtp_2 _14207_ (.CLK(clk),
    .D(_02836_),
    .Q(\data_array.data0[2][55] ));
 sky130_fd_sc_hd__dfxtp_2 _14208_ (.CLK(clk),
    .D(_02837_),
    .Q(\data_array.data0[2][56] ));
 sky130_fd_sc_hd__dfxtp_2 _14209_ (.CLK(clk),
    .D(_02838_),
    .Q(\data_array.data0[2][57] ));
 sky130_fd_sc_hd__dfxtp_2 _14210_ (.CLK(clk),
    .D(_02839_),
    .Q(\data_array.data0[2][58] ));
 sky130_fd_sc_hd__dfxtp_2 _14211_ (.CLK(clk),
    .D(_02840_),
    .Q(\data_array.data0[2][59] ));
 sky130_fd_sc_hd__dfxtp_2 _14212_ (.CLK(clk),
    .D(_02841_),
    .Q(\data_array.data0[2][60] ));
 sky130_fd_sc_hd__dfxtp_2 _14213_ (.CLK(clk),
    .D(_02842_),
    .Q(\data_array.data0[2][61] ));
 sky130_fd_sc_hd__dfxtp_2 _14214_ (.CLK(clk),
    .D(_02843_),
    .Q(\data_array.data0[2][62] ));
 sky130_fd_sc_hd__dfxtp_2 _14215_ (.CLK(clk),
    .D(_02844_),
    .Q(\data_array.data0[2][63] ));
 sky130_fd_sc_hd__dfxtp_2 _14216_ (.CLK(clk),
    .D(_02845_),
    .Q(\data_array.data1[12][0] ));
 sky130_fd_sc_hd__dfxtp_2 _14217_ (.CLK(clk),
    .D(_02846_),
    .Q(\data_array.data1[12][1] ));
 sky130_fd_sc_hd__dfxtp_2 _14218_ (.CLK(clk),
    .D(_02847_),
    .Q(\data_array.data1[12][2] ));
 sky130_fd_sc_hd__dfxtp_2 _14219_ (.CLK(clk),
    .D(_02848_),
    .Q(\data_array.data1[12][3] ));
 sky130_fd_sc_hd__dfxtp_2 _14220_ (.CLK(clk),
    .D(_02849_),
    .Q(\data_array.data1[12][4] ));
 sky130_fd_sc_hd__dfxtp_2 _14221_ (.CLK(clk),
    .D(_02850_),
    .Q(\data_array.data1[12][5] ));
 sky130_fd_sc_hd__dfxtp_2 _14222_ (.CLK(clk),
    .D(_02851_),
    .Q(\data_array.data1[12][6] ));
 sky130_fd_sc_hd__dfxtp_2 _14223_ (.CLK(clk),
    .D(_02852_),
    .Q(\data_array.data1[12][7] ));
 sky130_fd_sc_hd__dfxtp_2 _14224_ (.CLK(clk),
    .D(_02853_),
    .Q(\data_array.data1[12][8] ));
 sky130_fd_sc_hd__dfxtp_2 _14225_ (.CLK(clk),
    .D(_02854_),
    .Q(\data_array.data1[12][9] ));
 sky130_fd_sc_hd__dfxtp_2 _14226_ (.CLK(clk),
    .D(_02855_),
    .Q(\data_array.data1[12][10] ));
 sky130_fd_sc_hd__dfxtp_2 _14227_ (.CLK(clk),
    .D(_02856_),
    .Q(\data_array.data1[12][11] ));
 sky130_fd_sc_hd__dfxtp_2 _14228_ (.CLK(clk),
    .D(_02857_),
    .Q(\data_array.data1[12][12] ));
 sky130_fd_sc_hd__dfxtp_2 _14229_ (.CLK(clk),
    .D(_02858_),
    .Q(\data_array.data1[12][13] ));
 sky130_fd_sc_hd__dfxtp_2 _14230_ (.CLK(clk),
    .D(_02859_),
    .Q(\data_array.data1[12][14] ));
 sky130_fd_sc_hd__dfxtp_2 _14231_ (.CLK(clk),
    .D(_02860_),
    .Q(\data_array.data1[12][15] ));
 sky130_fd_sc_hd__dfxtp_2 _14232_ (.CLK(clk),
    .D(_02861_),
    .Q(\data_array.data1[12][16] ));
 sky130_fd_sc_hd__dfxtp_2 _14233_ (.CLK(clk),
    .D(_02862_),
    .Q(\data_array.data1[12][17] ));
 sky130_fd_sc_hd__dfxtp_2 _14234_ (.CLK(clk),
    .D(_02863_),
    .Q(\data_array.data1[12][18] ));
 sky130_fd_sc_hd__dfxtp_2 _14235_ (.CLK(clk),
    .D(_02864_),
    .Q(\data_array.data1[12][19] ));
 sky130_fd_sc_hd__dfxtp_2 _14236_ (.CLK(clk),
    .D(_02865_),
    .Q(\data_array.data1[12][20] ));
 sky130_fd_sc_hd__dfxtp_2 _14237_ (.CLK(clk),
    .D(_02866_),
    .Q(\data_array.data1[12][21] ));
 sky130_fd_sc_hd__dfxtp_2 _14238_ (.CLK(clk),
    .D(_02867_),
    .Q(\data_array.data1[12][22] ));
 sky130_fd_sc_hd__dfxtp_2 _14239_ (.CLK(clk),
    .D(_02868_),
    .Q(\data_array.data1[12][23] ));
 sky130_fd_sc_hd__dfxtp_2 _14240_ (.CLK(clk),
    .D(_02869_),
    .Q(\data_array.data1[12][24] ));
 sky130_fd_sc_hd__dfxtp_2 _14241_ (.CLK(clk),
    .D(_02870_),
    .Q(\data_array.data1[12][25] ));
 sky130_fd_sc_hd__dfxtp_2 _14242_ (.CLK(clk),
    .D(_02871_),
    .Q(\data_array.data1[12][26] ));
 sky130_fd_sc_hd__dfxtp_2 _14243_ (.CLK(clk),
    .D(_02872_),
    .Q(\data_array.data1[12][27] ));
 sky130_fd_sc_hd__dfxtp_2 _14244_ (.CLK(clk),
    .D(_02873_),
    .Q(\data_array.data1[12][28] ));
 sky130_fd_sc_hd__dfxtp_2 _14245_ (.CLK(clk),
    .D(_02874_),
    .Q(\data_array.data1[12][29] ));
 sky130_fd_sc_hd__dfxtp_2 _14246_ (.CLK(clk),
    .D(_02875_),
    .Q(\data_array.data1[12][30] ));
 sky130_fd_sc_hd__dfxtp_2 _14247_ (.CLK(clk),
    .D(_02876_),
    .Q(\data_array.data1[12][31] ));
 sky130_fd_sc_hd__dfxtp_2 _14248_ (.CLK(clk),
    .D(_02877_),
    .Q(\data_array.data1[12][32] ));
 sky130_fd_sc_hd__dfxtp_2 _14249_ (.CLK(clk),
    .D(_02878_),
    .Q(\data_array.data1[12][33] ));
 sky130_fd_sc_hd__dfxtp_2 _14250_ (.CLK(clk),
    .D(_02879_),
    .Q(\data_array.data1[12][34] ));
 sky130_fd_sc_hd__dfxtp_2 _14251_ (.CLK(clk),
    .D(_02880_),
    .Q(\data_array.data1[12][35] ));
 sky130_fd_sc_hd__dfxtp_2 _14252_ (.CLK(clk),
    .D(_02881_),
    .Q(\data_array.data1[12][36] ));
 sky130_fd_sc_hd__dfxtp_2 _14253_ (.CLK(clk),
    .D(_02882_),
    .Q(\data_array.data1[12][37] ));
 sky130_fd_sc_hd__dfxtp_2 _14254_ (.CLK(clk),
    .D(_02883_),
    .Q(\data_array.data1[12][38] ));
 sky130_fd_sc_hd__dfxtp_2 _14255_ (.CLK(clk),
    .D(_02884_),
    .Q(\data_array.data1[12][39] ));
 sky130_fd_sc_hd__dfxtp_2 _14256_ (.CLK(clk),
    .D(_02885_),
    .Q(\data_array.data1[12][40] ));
 sky130_fd_sc_hd__dfxtp_2 _14257_ (.CLK(clk),
    .D(_02886_),
    .Q(\data_array.data1[12][41] ));
 sky130_fd_sc_hd__dfxtp_2 _14258_ (.CLK(clk),
    .D(_02887_),
    .Q(\data_array.data1[12][42] ));
 sky130_fd_sc_hd__dfxtp_2 _14259_ (.CLK(clk),
    .D(_02888_),
    .Q(\data_array.data1[12][43] ));
 sky130_fd_sc_hd__dfxtp_2 _14260_ (.CLK(clk),
    .D(_02889_),
    .Q(\data_array.data1[12][44] ));
 sky130_fd_sc_hd__dfxtp_2 _14261_ (.CLK(clk),
    .D(_02890_),
    .Q(\data_array.data1[12][45] ));
 sky130_fd_sc_hd__dfxtp_2 _14262_ (.CLK(clk),
    .D(_02891_),
    .Q(\data_array.data1[12][46] ));
 sky130_fd_sc_hd__dfxtp_2 _14263_ (.CLK(clk),
    .D(_02892_),
    .Q(\data_array.data1[12][47] ));
 sky130_fd_sc_hd__dfxtp_2 _14264_ (.CLK(clk),
    .D(_02893_),
    .Q(\data_array.data1[12][48] ));
 sky130_fd_sc_hd__dfxtp_2 _14265_ (.CLK(clk),
    .D(_02894_),
    .Q(\data_array.data1[12][49] ));
 sky130_fd_sc_hd__dfxtp_2 _14266_ (.CLK(clk),
    .D(_02895_),
    .Q(\data_array.data1[12][50] ));
 sky130_fd_sc_hd__dfxtp_2 _14267_ (.CLK(clk),
    .D(_02896_),
    .Q(\data_array.data1[12][51] ));
 sky130_fd_sc_hd__dfxtp_2 _14268_ (.CLK(clk),
    .D(_02897_),
    .Q(\data_array.data1[12][52] ));
 sky130_fd_sc_hd__dfxtp_2 _14269_ (.CLK(clk),
    .D(_02898_),
    .Q(\data_array.data1[12][53] ));
 sky130_fd_sc_hd__dfxtp_2 _14270_ (.CLK(clk),
    .D(_02899_),
    .Q(\data_array.data1[12][54] ));
 sky130_fd_sc_hd__dfxtp_2 _14271_ (.CLK(clk),
    .D(_02900_),
    .Q(\data_array.data1[12][55] ));
 sky130_fd_sc_hd__dfxtp_2 _14272_ (.CLK(clk),
    .D(_02901_),
    .Q(\data_array.data1[12][56] ));
 sky130_fd_sc_hd__dfxtp_2 _14273_ (.CLK(clk),
    .D(_02902_),
    .Q(\data_array.data1[12][57] ));
 sky130_fd_sc_hd__dfxtp_2 _14274_ (.CLK(clk),
    .D(_02903_),
    .Q(\data_array.data1[12][58] ));
 sky130_fd_sc_hd__dfxtp_2 _14275_ (.CLK(clk),
    .D(_02904_),
    .Q(\data_array.data1[12][59] ));
 sky130_fd_sc_hd__dfxtp_2 _14276_ (.CLK(clk),
    .D(_02905_),
    .Q(\data_array.data1[12][60] ));
 sky130_fd_sc_hd__dfxtp_2 _14277_ (.CLK(clk),
    .D(_02906_),
    .Q(\data_array.data1[12][61] ));
 sky130_fd_sc_hd__dfxtp_2 _14278_ (.CLK(clk),
    .D(_02907_),
    .Q(\data_array.data1[12][62] ));
 sky130_fd_sc_hd__dfxtp_2 _14279_ (.CLK(clk),
    .D(_02908_),
    .Q(\data_array.data1[12][63] ));
 sky130_fd_sc_hd__dfxtp_2 _14280_ (.CLK(clk),
    .D(_02909_),
    .Q(\data_array.data1[11][0] ));
 sky130_fd_sc_hd__dfxtp_2 _14281_ (.CLK(clk),
    .D(_02910_),
    .Q(\data_array.data1[11][1] ));
 sky130_fd_sc_hd__dfxtp_2 _14282_ (.CLK(clk),
    .D(_02911_),
    .Q(\data_array.data1[11][2] ));
 sky130_fd_sc_hd__dfxtp_2 _14283_ (.CLK(clk),
    .D(_02912_),
    .Q(\data_array.data1[11][3] ));
 sky130_fd_sc_hd__dfxtp_2 _14284_ (.CLK(clk),
    .D(_02913_),
    .Q(\data_array.data1[11][4] ));
 sky130_fd_sc_hd__dfxtp_2 _14285_ (.CLK(clk),
    .D(_02914_),
    .Q(\data_array.data1[11][5] ));
 sky130_fd_sc_hd__dfxtp_2 _14286_ (.CLK(clk),
    .D(_02915_),
    .Q(\data_array.data1[11][6] ));
 sky130_fd_sc_hd__dfxtp_2 _14287_ (.CLK(clk),
    .D(_02916_),
    .Q(\data_array.data1[11][7] ));
 sky130_fd_sc_hd__dfxtp_2 _14288_ (.CLK(clk),
    .D(_02917_),
    .Q(\data_array.data1[11][8] ));
 sky130_fd_sc_hd__dfxtp_2 _14289_ (.CLK(clk),
    .D(_02918_),
    .Q(\data_array.data1[11][9] ));
 sky130_fd_sc_hd__dfxtp_2 _14290_ (.CLK(clk),
    .D(_02919_),
    .Q(\data_array.data1[11][10] ));
 sky130_fd_sc_hd__dfxtp_2 _14291_ (.CLK(clk),
    .D(_02920_),
    .Q(\data_array.data1[11][11] ));
 sky130_fd_sc_hd__dfxtp_2 _14292_ (.CLK(clk),
    .D(_02921_),
    .Q(\data_array.data1[11][12] ));
 sky130_fd_sc_hd__dfxtp_2 _14293_ (.CLK(clk),
    .D(_02922_),
    .Q(\data_array.data1[11][13] ));
 sky130_fd_sc_hd__dfxtp_2 _14294_ (.CLK(clk),
    .D(_02923_),
    .Q(\data_array.data1[11][14] ));
 sky130_fd_sc_hd__dfxtp_2 _14295_ (.CLK(clk),
    .D(_02924_),
    .Q(\data_array.data1[11][15] ));
 sky130_fd_sc_hd__dfxtp_2 _14296_ (.CLK(clk),
    .D(_02925_),
    .Q(\data_array.data1[11][16] ));
 sky130_fd_sc_hd__dfxtp_2 _14297_ (.CLK(clk),
    .D(_02926_),
    .Q(\data_array.data1[11][17] ));
 sky130_fd_sc_hd__dfxtp_2 _14298_ (.CLK(clk),
    .D(_02927_),
    .Q(\data_array.data1[11][18] ));
 sky130_fd_sc_hd__dfxtp_2 _14299_ (.CLK(clk),
    .D(_02928_),
    .Q(\data_array.data1[11][19] ));
 sky130_fd_sc_hd__dfxtp_2 _14300_ (.CLK(clk),
    .D(_02929_),
    .Q(\data_array.data1[11][20] ));
 sky130_fd_sc_hd__dfxtp_2 _14301_ (.CLK(clk),
    .D(_02930_),
    .Q(\data_array.data1[11][21] ));
 sky130_fd_sc_hd__dfxtp_2 _14302_ (.CLK(clk),
    .D(_02931_),
    .Q(\data_array.data1[11][22] ));
 sky130_fd_sc_hd__dfxtp_2 _14303_ (.CLK(clk),
    .D(_02932_),
    .Q(\data_array.data1[11][23] ));
 sky130_fd_sc_hd__dfxtp_2 _14304_ (.CLK(clk),
    .D(_02933_),
    .Q(\data_array.data1[11][24] ));
 sky130_fd_sc_hd__dfxtp_2 _14305_ (.CLK(clk),
    .D(_02934_),
    .Q(\data_array.data1[11][25] ));
 sky130_fd_sc_hd__dfxtp_2 _14306_ (.CLK(clk),
    .D(_02935_),
    .Q(\data_array.data1[11][26] ));
 sky130_fd_sc_hd__dfxtp_2 _14307_ (.CLK(clk),
    .D(_02936_),
    .Q(\data_array.data1[11][27] ));
 sky130_fd_sc_hd__dfxtp_2 _14308_ (.CLK(clk),
    .D(_02937_),
    .Q(\data_array.data1[11][28] ));
 sky130_fd_sc_hd__dfxtp_2 _14309_ (.CLK(clk),
    .D(_02938_),
    .Q(\data_array.data1[11][29] ));
 sky130_fd_sc_hd__dfxtp_2 _14310_ (.CLK(clk),
    .D(_02939_),
    .Q(\data_array.data1[11][30] ));
 sky130_fd_sc_hd__dfxtp_2 _14311_ (.CLK(clk),
    .D(_02940_),
    .Q(\data_array.data1[11][31] ));
 sky130_fd_sc_hd__dfxtp_2 _14312_ (.CLK(clk),
    .D(_02941_),
    .Q(\data_array.data1[11][32] ));
 sky130_fd_sc_hd__dfxtp_2 _14313_ (.CLK(clk),
    .D(_02942_),
    .Q(\data_array.data1[11][33] ));
 sky130_fd_sc_hd__dfxtp_2 _14314_ (.CLK(clk),
    .D(_02943_),
    .Q(\data_array.data1[11][34] ));
 sky130_fd_sc_hd__dfxtp_2 _14315_ (.CLK(clk),
    .D(_02944_),
    .Q(\data_array.data1[11][35] ));
 sky130_fd_sc_hd__dfxtp_2 _14316_ (.CLK(clk),
    .D(_02945_),
    .Q(\data_array.data1[11][36] ));
 sky130_fd_sc_hd__dfxtp_2 _14317_ (.CLK(clk),
    .D(_02946_),
    .Q(\data_array.data1[11][37] ));
 sky130_fd_sc_hd__dfxtp_2 _14318_ (.CLK(clk),
    .D(_02947_),
    .Q(\data_array.data1[11][38] ));
 sky130_fd_sc_hd__dfxtp_2 _14319_ (.CLK(clk),
    .D(_02948_),
    .Q(\data_array.data1[11][39] ));
 sky130_fd_sc_hd__dfxtp_2 _14320_ (.CLK(clk),
    .D(_02949_),
    .Q(\data_array.data1[11][40] ));
 sky130_fd_sc_hd__dfxtp_2 _14321_ (.CLK(clk),
    .D(_02950_),
    .Q(\data_array.data1[11][41] ));
 sky130_fd_sc_hd__dfxtp_2 _14322_ (.CLK(clk),
    .D(_02951_),
    .Q(\data_array.data1[11][42] ));
 sky130_fd_sc_hd__dfxtp_2 _14323_ (.CLK(clk),
    .D(_02952_),
    .Q(\data_array.data1[11][43] ));
 sky130_fd_sc_hd__dfxtp_2 _14324_ (.CLK(clk),
    .D(_02953_),
    .Q(\data_array.data1[11][44] ));
 sky130_fd_sc_hd__dfxtp_2 _14325_ (.CLK(clk),
    .D(_02954_),
    .Q(\data_array.data1[11][45] ));
 sky130_fd_sc_hd__dfxtp_2 _14326_ (.CLK(clk),
    .D(_02955_),
    .Q(\data_array.data1[11][46] ));
 sky130_fd_sc_hd__dfxtp_2 _14327_ (.CLK(clk),
    .D(_02956_),
    .Q(\data_array.data1[11][47] ));
 sky130_fd_sc_hd__dfxtp_2 _14328_ (.CLK(clk),
    .D(_02957_),
    .Q(\data_array.data1[11][48] ));
 sky130_fd_sc_hd__dfxtp_2 _14329_ (.CLK(clk),
    .D(_02958_),
    .Q(\data_array.data1[11][49] ));
 sky130_fd_sc_hd__dfxtp_2 _14330_ (.CLK(clk),
    .D(_02959_),
    .Q(\data_array.data1[11][50] ));
 sky130_fd_sc_hd__dfxtp_2 _14331_ (.CLK(clk),
    .D(_02960_),
    .Q(\data_array.data1[11][51] ));
 sky130_fd_sc_hd__dfxtp_2 _14332_ (.CLK(clk),
    .D(_02961_),
    .Q(\data_array.data1[11][52] ));
 sky130_fd_sc_hd__dfxtp_2 _14333_ (.CLK(clk),
    .D(_02962_),
    .Q(\data_array.data1[11][53] ));
 sky130_fd_sc_hd__dfxtp_2 _14334_ (.CLK(clk),
    .D(_02963_),
    .Q(\data_array.data1[11][54] ));
 sky130_fd_sc_hd__dfxtp_2 _14335_ (.CLK(clk),
    .D(_02964_),
    .Q(\data_array.data1[11][55] ));
 sky130_fd_sc_hd__dfxtp_2 _14336_ (.CLK(clk),
    .D(_02965_),
    .Q(\data_array.data1[11][56] ));
 sky130_fd_sc_hd__dfxtp_2 _14337_ (.CLK(clk),
    .D(_02966_),
    .Q(\data_array.data1[11][57] ));
 sky130_fd_sc_hd__dfxtp_2 _14338_ (.CLK(clk),
    .D(_02967_),
    .Q(\data_array.data1[11][58] ));
 sky130_fd_sc_hd__dfxtp_2 _14339_ (.CLK(clk),
    .D(_02968_),
    .Q(\data_array.data1[11][59] ));
 sky130_fd_sc_hd__dfxtp_2 _14340_ (.CLK(clk),
    .D(_02969_),
    .Q(\data_array.data1[11][60] ));
 sky130_fd_sc_hd__dfxtp_2 _14341_ (.CLK(clk),
    .D(_02970_),
    .Q(\data_array.data1[11][61] ));
 sky130_fd_sc_hd__dfxtp_2 _14342_ (.CLK(clk),
    .D(_02971_),
    .Q(\data_array.data1[11][62] ));
 sky130_fd_sc_hd__dfxtp_2 _14343_ (.CLK(clk),
    .D(_02972_),
    .Q(\data_array.data1[11][63] ));
 sky130_fd_sc_hd__dfstp_2 _14344_ (.CLK(clk),
    .D(_00186_),
    .SET_B(_00189_),
    .Q(\fsm.state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _14345_ (.CLK(clk),
    .D(_00187_),
    .RESET_B(_00190_),
    .Q(mem_write));
 sky130_fd_sc_hd__dfrtp_2 _14346_ (.CLK(clk),
    .D(_00183_),
    .RESET_B(_00191_),
    .Q(\fsm.state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _14347_ (.CLK(clk),
    .D(_00184_),
    .RESET_B(_00192_),
    .Q(\fsm.state[3] ));
 sky130_fd_sc_hd__dfrtp_2 _14348_ (.CLK(clk),
    .D(_00188_),
    .RESET_B(_00193_),
    .Q(mem_read));
 sky130_fd_sc_hd__dfrtp_2 _14349_ (.CLK(clk),
    .D(_00185_),
    .RESET_B(_00194_),
    .Q(\fsm.state[5] ));
 sky130_fd_sc_hd__dfxtp_2 _14350_ (.CLK(clk),
    .D(_02973_),
    .Q(\data_array.data1[10][0] ));
 sky130_fd_sc_hd__dfxtp_2 _14351_ (.CLK(clk),
    .D(_02974_),
    .Q(\data_array.data1[10][1] ));
 sky130_fd_sc_hd__dfxtp_2 _14352_ (.CLK(clk),
    .D(_02975_),
    .Q(\data_array.data1[10][2] ));
 sky130_fd_sc_hd__dfxtp_2 _14353_ (.CLK(clk),
    .D(_02976_),
    .Q(\data_array.data1[10][3] ));
 sky130_fd_sc_hd__dfxtp_2 _14354_ (.CLK(clk),
    .D(_02977_),
    .Q(\data_array.data1[10][4] ));
 sky130_fd_sc_hd__dfxtp_2 _14355_ (.CLK(clk),
    .D(_02978_),
    .Q(\data_array.data1[10][5] ));
 sky130_fd_sc_hd__dfxtp_2 _14356_ (.CLK(clk),
    .D(_02979_),
    .Q(\data_array.data1[10][6] ));
 sky130_fd_sc_hd__dfxtp_2 _14357_ (.CLK(clk),
    .D(_02980_),
    .Q(\data_array.data1[10][7] ));
 sky130_fd_sc_hd__dfxtp_2 _14358_ (.CLK(clk),
    .D(_02981_),
    .Q(\data_array.data1[10][8] ));
 sky130_fd_sc_hd__dfxtp_2 _14359_ (.CLK(clk),
    .D(_02982_),
    .Q(\data_array.data1[10][9] ));
 sky130_fd_sc_hd__dfxtp_2 _14360_ (.CLK(clk),
    .D(_02983_),
    .Q(\data_array.data1[10][10] ));
 sky130_fd_sc_hd__dfxtp_2 _14361_ (.CLK(clk),
    .D(_02984_),
    .Q(\data_array.data1[10][11] ));
 sky130_fd_sc_hd__dfxtp_2 _14362_ (.CLK(clk),
    .D(_02985_),
    .Q(\data_array.data1[10][12] ));
 sky130_fd_sc_hd__dfxtp_2 _14363_ (.CLK(clk),
    .D(_02986_),
    .Q(\data_array.data1[10][13] ));
 sky130_fd_sc_hd__dfxtp_2 _14364_ (.CLK(clk),
    .D(_02987_),
    .Q(\data_array.data1[10][14] ));
 sky130_fd_sc_hd__dfxtp_2 _14365_ (.CLK(clk),
    .D(_02988_),
    .Q(\data_array.data1[10][15] ));
 sky130_fd_sc_hd__dfxtp_2 _14366_ (.CLK(clk),
    .D(_02989_),
    .Q(\data_array.data1[10][16] ));
 sky130_fd_sc_hd__dfxtp_2 _14367_ (.CLK(clk),
    .D(_02990_),
    .Q(\data_array.data1[10][17] ));
 sky130_fd_sc_hd__dfxtp_2 _14368_ (.CLK(clk),
    .D(_02991_),
    .Q(\data_array.data1[10][18] ));
 sky130_fd_sc_hd__dfxtp_2 _14369_ (.CLK(clk),
    .D(_02992_),
    .Q(\data_array.data1[10][19] ));
 sky130_fd_sc_hd__dfxtp_2 _14370_ (.CLK(clk),
    .D(_02993_),
    .Q(\data_array.data1[10][20] ));
 sky130_fd_sc_hd__dfxtp_2 _14371_ (.CLK(clk),
    .D(_02994_),
    .Q(\data_array.data1[10][21] ));
 sky130_fd_sc_hd__dfxtp_2 _14372_ (.CLK(clk),
    .D(_02995_),
    .Q(\data_array.data1[10][22] ));
 sky130_fd_sc_hd__dfxtp_2 _14373_ (.CLK(clk),
    .D(_02996_),
    .Q(\data_array.data1[10][23] ));
 sky130_fd_sc_hd__dfxtp_2 _14374_ (.CLK(clk),
    .D(_02997_),
    .Q(\data_array.data1[10][24] ));
 sky130_fd_sc_hd__dfxtp_2 _14375_ (.CLK(clk),
    .D(_02998_),
    .Q(\data_array.data1[10][25] ));
 sky130_fd_sc_hd__dfxtp_2 _14376_ (.CLK(clk),
    .D(_02999_),
    .Q(\data_array.data1[10][26] ));
 sky130_fd_sc_hd__dfxtp_2 _14377_ (.CLK(clk),
    .D(_03000_),
    .Q(\data_array.data1[10][27] ));
 sky130_fd_sc_hd__dfxtp_2 _14378_ (.CLK(clk),
    .D(_03001_),
    .Q(\data_array.data1[10][28] ));
 sky130_fd_sc_hd__dfxtp_2 _14379_ (.CLK(clk),
    .D(_03002_),
    .Q(\data_array.data1[10][29] ));
 sky130_fd_sc_hd__dfxtp_2 _14380_ (.CLK(clk),
    .D(_03003_),
    .Q(\data_array.data1[10][30] ));
 sky130_fd_sc_hd__dfxtp_2 _14381_ (.CLK(clk),
    .D(_03004_),
    .Q(\data_array.data1[10][31] ));
 sky130_fd_sc_hd__dfxtp_2 _14382_ (.CLK(clk),
    .D(_03005_),
    .Q(\data_array.data1[10][32] ));
 sky130_fd_sc_hd__dfxtp_2 _14383_ (.CLK(clk),
    .D(_03006_),
    .Q(\data_array.data1[10][33] ));
 sky130_fd_sc_hd__dfxtp_2 _14384_ (.CLK(clk),
    .D(_03007_),
    .Q(\data_array.data1[10][34] ));
 sky130_fd_sc_hd__dfxtp_2 _14385_ (.CLK(clk),
    .D(_03008_),
    .Q(\data_array.data1[10][35] ));
 sky130_fd_sc_hd__dfxtp_2 _14386_ (.CLK(clk),
    .D(_03009_),
    .Q(\data_array.data1[10][36] ));
 sky130_fd_sc_hd__dfxtp_2 _14387_ (.CLK(clk),
    .D(_03010_),
    .Q(\data_array.data1[10][37] ));
 sky130_fd_sc_hd__dfxtp_2 _14388_ (.CLK(clk),
    .D(_03011_),
    .Q(\data_array.data1[10][38] ));
 sky130_fd_sc_hd__dfxtp_2 _14389_ (.CLK(clk),
    .D(_03012_),
    .Q(\data_array.data1[10][39] ));
 sky130_fd_sc_hd__dfxtp_2 _14390_ (.CLK(clk),
    .D(_03013_),
    .Q(\data_array.data1[10][40] ));
 sky130_fd_sc_hd__dfxtp_2 _14391_ (.CLK(clk),
    .D(_03014_),
    .Q(\data_array.data1[10][41] ));
 sky130_fd_sc_hd__dfxtp_2 _14392_ (.CLK(clk),
    .D(_03015_),
    .Q(\data_array.data1[10][42] ));
 sky130_fd_sc_hd__dfxtp_2 _14393_ (.CLK(clk),
    .D(_03016_),
    .Q(\data_array.data1[10][43] ));
 sky130_fd_sc_hd__dfxtp_2 _14394_ (.CLK(clk),
    .D(_03017_),
    .Q(\data_array.data1[10][44] ));
 sky130_fd_sc_hd__dfxtp_2 _14395_ (.CLK(clk),
    .D(_03018_),
    .Q(\data_array.data1[10][45] ));
 sky130_fd_sc_hd__dfxtp_2 _14396_ (.CLK(clk),
    .D(_03019_),
    .Q(\data_array.data1[10][46] ));
 sky130_fd_sc_hd__dfxtp_2 _14397_ (.CLK(clk),
    .D(_03020_),
    .Q(\data_array.data1[10][47] ));
 sky130_fd_sc_hd__dfxtp_2 _14398_ (.CLK(clk),
    .D(_03021_),
    .Q(\data_array.data1[10][48] ));
 sky130_fd_sc_hd__dfxtp_2 _14399_ (.CLK(clk),
    .D(_03022_),
    .Q(\data_array.data1[10][49] ));
 sky130_fd_sc_hd__dfxtp_2 _14400_ (.CLK(clk),
    .D(_03023_),
    .Q(\data_array.data1[10][50] ));
 sky130_fd_sc_hd__dfxtp_2 _14401_ (.CLK(clk),
    .D(_03024_),
    .Q(\data_array.data1[10][51] ));
 sky130_fd_sc_hd__dfxtp_2 _14402_ (.CLK(clk),
    .D(_03025_),
    .Q(\data_array.data1[10][52] ));
 sky130_fd_sc_hd__dfxtp_2 _14403_ (.CLK(clk),
    .D(_03026_),
    .Q(\data_array.data1[10][53] ));
 sky130_fd_sc_hd__dfxtp_2 _14404_ (.CLK(clk),
    .D(_03027_),
    .Q(\data_array.data1[10][54] ));
 sky130_fd_sc_hd__dfxtp_2 _14405_ (.CLK(clk),
    .D(_03028_),
    .Q(\data_array.data1[10][55] ));
 sky130_fd_sc_hd__dfxtp_2 _14406_ (.CLK(clk),
    .D(_03029_),
    .Q(\data_array.data1[10][56] ));
 sky130_fd_sc_hd__dfxtp_2 _14407_ (.CLK(clk),
    .D(_03030_),
    .Q(\data_array.data1[10][57] ));
 sky130_fd_sc_hd__dfxtp_2 _14408_ (.CLK(clk),
    .D(_03031_),
    .Q(\data_array.data1[10][58] ));
 sky130_fd_sc_hd__dfxtp_2 _14409_ (.CLK(clk),
    .D(_03032_),
    .Q(\data_array.data1[10][59] ));
 sky130_fd_sc_hd__dfxtp_2 _14410_ (.CLK(clk),
    .D(_03033_),
    .Q(\data_array.data1[10][60] ));
 sky130_fd_sc_hd__dfxtp_2 _14411_ (.CLK(clk),
    .D(_03034_),
    .Q(\data_array.data1[10][61] ));
 sky130_fd_sc_hd__dfxtp_2 _14412_ (.CLK(clk),
    .D(_03035_),
    .Q(\data_array.data1[10][62] ));
 sky130_fd_sc_hd__dfxtp_2 _14413_ (.CLK(clk),
    .D(_03036_),
    .Q(\data_array.data1[10][63] ));
 sky130_fd_sc_hd__dfxtp_2 _14414_ (.CLK(clk),
    .D(_03037_),
    .Q(\lru_array.lru_mem[13] ));
 sky130_fd_sc_hd__dfxtp_2 _14415_ (.CLK(clk),
    .D(_03038_),
    .Q(\lru_array.lru_mem[14] ));
 sky130_fd_sc_hd__dfxtp_2 _14416_ (.CLK(clk),
    .D(_03039_),
    .Q(\data_array.data1[7][0] ));
 sky130_fd_sc_hd__dfxtp_2 _14417_ (.CLK(clk),
    .D(_03040_),
    .Q(\data_array.data1[7][1] ));
 sky130_fd_sc_hd__dfxtp_2 _14418_ (.CLK(clk),
    .D(_03041_),
    .Q(\data_array.data1[7][2] ));
 sky130_fd_sc_hd__dfxtp_2 _14419_ (.CLK(clk),
    .D(_03042_),
    .Q(\data_array.data1[7][3] ));
 sky130_fd_sc_hd__dfxtp_2 _14420_ (.CLK(clk),
    .D(_03043_),
    .Q(\data_array.data1[7][4] ));
 sky130_fd_sc_hd__dfxtp_2 _14421_ (.CLK(clk),
    .D(_03044_),
    .Q(\data_array.data1[7][5] ));
 sky130_fd_sc_hd__dfxtp_2 _14422_ (.CLK(clk),
    .D(_03045_),
    .Q(\data_array.data1[7][6] ));
 sky130_fd_sc_hd__dfxtp_2 _14423_ (.CLK(clk),
    .D(_03046_),
    .Q(\data_array.data1[7][7] ));
 sky130_fd_sc_hd__dfxtp_2 _14424_ (.CLK(clk),
    .D(_03047_),
    .Q(\data_array.data1[7][8] ));
 sky130_fd_sc_hd__dfxtp_2 _14425_ (.CLK(clk),
    .D(_03048_),
    .Q(\data_array.data1[7][9] ));
 sky130_fd_sc_hd__dfxtp_2 _14426_ (.CLK(clk),
    .D(_03049_),
    .Q(\data_array.data1[7][10] ));
 sky130_fd_sc_hd__dfxtp_2 _14427_ (.CLK(clk),
    .D(_03050_),
    .Q(\data_array.data1[7][11] ));
 sky130_fd_sc_hd__dfxtp_2 _14428_ (.CLK(clk),
    .D(_03051_),
    .Q(\data_array.data1[7][12] ));
 sky130_fd_sc_hd__dfxtp_2 _14429_ (.CLK(clk),
    .D(_03052_),
    .Q(\data_array.data1[7][13] ));
 sky130_fd_sc_hd__dfxtp_2 _14430_ (.CLK(clk),
    .D(_03053_),
    .Q(\data_array.data1[7][14] ));
 sky130_fd_sc_hd__dfxtp_2 _14431_ (.CLK(clk),
    .D(_03054_),
    .Q(\data_array.data1[7][15] ));
 sky130_fd_sc_hd__dfxtp_2 _14432_ (.CLK(clk),
    .D(_03055_),
    .Q(\data_array.data1[7][16] ));
 sky130_fd_sc_hd__dfxtp_2 _14433_ (.CLK(clk),
    .D(_03056_),
    .Q(\data_array.data1[7][17] ));
 sky130_fd_sc_hd__dfxtp_2 _14434_ (.CLK(clk),
    .D(_03057_),
    .Q(\data_array.data1[7][18] ));
 sky130_fd_sc_hd__dfxtp_2 _14435_ (.CLK(clk),
    .D(_03058_),
    .Q(\data_array.data1[7][19] ));
 sky130_fd_sc_hd__dfxtp_2 _14436_ (.CLK(clk),
    .D(_03059_),
    .Q(\data_array.data1[7][20] ));
 sky130_fd_sc_hd__dfxtp_2 _14437_ (.CLK(clk),
    .D(_03060_),
    .Q(\data_array.data1[7][21] ));
 sky130_fd_sc_hd__dfxtp_2 _14438_ (.CLK(clk),
    .D(_03061_),
    .Q(\data_array.data1[7][22] ));
 sky130_fd_sc_hd__dfxtp_2 _14439_ (.CLK(clk),
    .D(_03062_),
    .Q(\data_array.data1[7][23] ));
 sky130_fd_sc_hd__dfxtp_2 _14440_ (.CLK(clk),
    .D(_03063_),
    .Q(\data_array.data1[7][24] ));
 sky130_fd_sc_hd__dfxtp_2 _14441_ (.CLK(clk),
    .D(_03064_),
    .Q(\data_array.data1[7][25] ));
 sky130_fd_sc_hd__dfxtp_2 _14442_ (.CLK(clk),
    .D(_03065_),
    .Q(\data_array.data1[7][26] ));
 sky130_fd_sc_hd__dfxtp_2 _14443_ (.CLK(clk),
    .D(_03066_),
    .Q(\data_array.data1[7][27] ));
 sky130_fd_sc_hd__dfxtp_2 _14444_ (.CLK(clk),
    .D(_03067_),
    .Q(\data_array.data1[7][28] ));
 sky130_fd_sc_hd__dfxtp_2 _14445_ (.CLK(clk),
    .D(_03068_),
    .Q(\data_array.data1[7][29] ));
 sky130_fd_sc_hd__dfxtp_2 _14446_ (.CLK(clk),
    .D(_03069_),
    .Q(\data_array.data1[7][30] ));
 sky130_fd_sc_hd__dfxtp_2 _14447_ (.CLK(clk),
    .D(_03070_),
    .Q(\data_array.data1[7][31] ));
 sky130_fd_sc_hd__dfxtp_2 _14448_ (.CLK(clk),
    .D(_03071_),
    .Q(\data_array.data1[7][32] ));
 sky130_fd_sc_hd__dfxtp_2 _14449_ (.CLK(clk),
    .D(_03072_),
    .Q(\data_array.data1[7][33] ));
 sky130_fd_sc_hd__dfxtp_2 _14450_ (.CLK(clk),
    .D(_03073_),
    .Q(\data_array.data1[7][34] ));
 sky130_fd_sc_hd__dfxtp_2 _14451_ (.CLK(clk),
    .D(_03074_),
    .Q(\data_array.data1[7][35] ));
 sky130_fd_sc_hd__dfxtp_2 _14452_ (.CLK(clk),
    .D(_03075_),
    .Q(\data_array.data1[7][36] ));
 sky130_fd_sc_hd__dfxtp_2 _14453_ (.CLK(clk),
    .D(_03076_),
    .Q(\data_array.data1[7][37] ));
 sky130_fd_sc_hd__dfxtp_2 _14454_ (.CLK(clk),
    .D(_03077_),
    .Q(\data_array.data1[7][38] ));
 sky130_fd_sc_hd__dfxtp_2 _14455_ (.CLK(clk),
    .D(_03078_),
    .Q(\data_array.data1[7][39] ));
 sky130_fd_sc_hd__dfxtp_2 _14456_ (.CLK(clk),
    .D(_03079_),
    .Q(\data_array.data1[7][40] ));
 sky130_fd_sc_hd__dfxtp_2 _14457_ (.CLK(clk),
    .D(_03080_),
    .Q(\data_array.data1[7][41] ));
 sky130_fd_sc_hd__dfxtp_2 _14458_ (.CLK(clk),
    .D(_03081_),
    .Q(\data_array.data1[7][42] ));
 sky130_fd_sc_hd__dfxtp_2 _14459_ (.CLK(clk),
    .D(_03082_),
    .Q(\data_array.data1[7][43] ));
 sky130_fd_sc_hd__dfxtp_2 _14460_ (.CLK(clk),
    .D(_03083_),
    .Q(\data_array.data1[7][44] ));
 sky130_fd_sc_hd__dfxtp_2 _14461_ (.CLK(clk),
    .D(_03084_),
    .Q(\data_array.data1[7][45] ));
 sky130_fd_sc_hd__dfxtp_2 _14462_ (.CLK(clk),
    .D(_03085_),
    .Q(\data_array.data1[7][46] ));
 sky130_fd_sc_hd__dfxtp_2 _14463_ (.CLK(clk),
    .D(_03086_),
    .Q(\data_array.data1[7][47] ));
 sky130_fd_sc_hd__dfxtp_2 _14464_ (.CLK(clk),
    .D(_03087_),
    .Q(\data_array.data1[7][48] ));
 sky130_fd_sc_hd__dfxtp_2 _14465_ (.CLK(clk),
    .D(_03088_),
    .Q(\data_array.data1[7][49] ));
 sky130_fd_sc_hd__dfxtp_2 _14466_ (.CLK(clk),
    .D(_03089_),
    .Q(\data_array.data1[7][50] ));
 sky130_fd_sc_hd__dfxtp_2 _14467_ (.CLK(clk),
    .D(_03090_),
    .Q(\data_array.data1[7][51] ));
 sky130_fd_sc_hd__dfxtp_2 _14468_ (.CLK(clk),
    .D(_03091_),
    .Q(\data_array.data1[7][52] ));
 sky130_fd_sc_hd__dfxtp_2 _14469_ (.CLK(clk),
    .D(_03092_),
    .Q(\data_array.data1[7][53] ));
 sky130_fd_sc_hd__dfxtp_2 _14470_ (.CLK(clk),
    .D(_03093_),
    .Q(\data_array.data1[7][54] ));
 sky130_fd_sc_hd__dfxtp_2 _14471_ (.CLK(clk),
    .D(_03094_),
    .Q(\data_array.data1[7][55] ));
 sky130_fd_sc_hd__dfxtp_2 _14472_ (.CLK(clk),
    .D(_03095_),
    .Q(\data_array.data1[7][56] ));
 sky130_fd_sc_hd__dfxtp_2 _14473_ (.CLK(clk),
    .D(_03096_),
    .Q(\data_array.data1[7][57] ));
 sky130_fd_sc_hd__dfxtp_2 _14474_ (.CLK(clk),
    .D(_03097_),
    .Q(\data_array.data1[7][58] ));
 sky130_fd_sc_hd__dfxtp_2 _14475_ (.CLK(clk),
    .D(_03098_),
    .Q(\data_array.data1[7][59] ));
 sky130_fd_sc_hd__dfxtp_2 _14476_ (.CLK(clk),
    .D(_03099_),
    .Q(\data_array.data1[7][60] ));
 sky130_fd_sc_hd__dfxtp_2 _14477_ (.CLK(clk),
    .D(_03100_),
    .Q(\data_array.data1[7][61] ));
 sky130_fd_sc_hd__dfxtp_2 _14478_ (.CLK(clk),
    .D(_03101_),
    .Q(\data_array.data1[7][62] ));
 sky130_fd_sc_hd__dfxtp_2 _14479_ (.CLK(clk),
    .D(_03102_),
    .Q(\data_array.data1[7][63] ));
 sky130_fd_sc_hd__dfxtp_2 _14480_ (.CLK(clk),
    .D(_03103_),
    .Q(\lru_array.lru_mem[9] ));
 sky130_fd_sc_hd__dfxtp_2 _14481_ (.CLK(clk),
    .D(_03104_),
    .Q(\tag_array.dirty0[15] ));
 sky130_fd_sc_hd__dfxtp_2 _14482_ (.CLK(clk),
    .D(_03105_),
    .Q(\tag_array.dirty0[1] ));
 sky130_fd_sc_hd__dfxtp_2 _14483_ (.CLK(clk),
    .D(_03106_),
    .Q(\tag_array.dirty0[2] ));
 sky130_fd_sc_hd__dfxtp_2 _14484_ (.CLK(clk),
    .D(_03107_),
    .Q(\tag_array.dirty0[3] ));
 sky130_fd_sc_hd__dfxtp_2 _14485_ (.CLK(clk),
    .D(_03108_),
    .Q(\tag_array.dirty0[4] ));
 sky130_fd_sc_hd__dfxtp_2 _14486_ (.CLK(clk),
    .D(_03109_),
    .Q(\tag_array.dirty0[5] ));
 sky130_fd_sc_hd__dfxtp_2 _14487_ (.CLK(clk),
    .D(_03110_),
    .Q(\tag_array.dirty0[6] ));
 sky130_fd_sc_hd__dfxtp_2 _14488_ (.CLK(clk),
    .D(_03111_),
    .Q(\tag_array.dirty0[7] ));
 sky130_fd_sc_hd__dfxtp_2 _14489_ (.CLK(clk),
    .D(_03112_),
    .Q(\tag_array.dirty0[8] ));
 sky130_fd_sc_hd__dfxtp_2 _14490_ (.CLK(clk),
    .D(_03113_),
    .Q(\tag_array.dirty0[0] ));
 sky130_fd_sc_hd__dfxtp_2 _14491_ (.CLK(clk),
    .D(_03114_),
    .Q(\tag_array.dirty0[10] ));
 sky130_fd_sc_hd__dfxtp_2 _14492_ (.CLK(clk),
    .D(_03115_),
    .Q(\tag_array.dirty0[11] ));
 sky130_fd_sc_hd__dfxtp_2 _14493_ (.CLK(clk),
    .D(_03116_),
    .Q(\tag_array.dirty0[12] ));
 sky130_fd_sc_hd__dfxtp_2 _14494_ (.CLK(clk),
    .D(_03117_),
    .Q(\tag_array.dirty0[13] ));
 sky130_fd_sc_hd__dfxtp_2 _14495_ (.CLK(clk),
    .D(_03118_),
    .Q(\lru_array.lru_mem[3] ));
 sky130_fd_sc_hd__dfxtp_2 _14496_ (.CLK(clk),
    .D(_03119_),
    .Q(\tag_array.dirty0[14] ));
 sky130_fd_sc_hd__dfxtp_2 _14497_ (.CLK(clk),
    .D(_00129_),
    .Q(dirty_way0));
 sky130_fd_sc_hd__dfxtp_2 _14498_ (.CLK(clk),
    .D(_03120_),
    .Q(\lru_array.lru_mem[12] ));
 sky130_fd_sc_hd__dfxtp_2 _14499_ (.CLK(clk),
    .D(_00128_),
    .Q(\fsm.lru_out ));
 sky130_fd_sc_hd__dfxtp_2 _14500_ (.CLK(clk),
    .D(_03121_),
    .Q(\lru_array.lru_mem[4] ));
 sky130_fd_sc_hd__dfxtp_2 _14501_ (.CLK(clk),
    .D(_03122_),
    .Q(\lru_array.lru_mem[5] ));
endmodule
